module pagerank_tb;

localparam N=64;
localparam WIDTH=16; //PLEASE UPDATE AS REQUIRED

reg clk; 
reg reset; 
always begin 
  #1 clk  = 1; 
  #1 clk = 0; 
end 

reg [N*N-1:0] adj; 
reg [N*WIDTH-1:0] nodeWeight; 

wire [10*WIDTH-1:0] top10Vals; 
wire [10*6-1:0] top10IDs; //N = 64, so at most 6 bits required

wire [WIDTH-1:0] nodeVal0; 
 wire [WIDTH-1:0] nodeVal16; 
 wire [WIDTH-1:0] nodeVal32; 
 wire [WIDTH-1:0] nodeVal48; 
pageRank #(N,WIDTH) pr(clk,reset,adj,nodeWeight,top10Vals,top10IDs,nodeVal0,nodeVal16,nodeVal32,nodeVal48);//PLEASE UPDATE AS PER YOUR MODULE DEFN

integer i; 

initial begin 
  reset = 0; 
  #1 reset = 1; 

for(i=0;i<N*N;i=i+1)begin 
  adj[i]=0; 
 end 
  adj[1] = 1; 
  adj[29] = 1; 
  adj[63] = 1; 
  adj[64] = 1; 
  adj[66] = 1; 
  adj[129] = 1; 
  adj[131] = 1; 
  adj[141] = 1; 
  adj[194] = 1; 
  adj[196] = 1; 
  adj[208] = 1; 
  adj[259] = 1; 
  adj[261] = 1; 
  adj[269] = 1; 
  adj[324] = 1; 
  adj[326] = 1; 
  adj[364] = 1; 
  adj[389] = 1; 
  adj[391] = 1; 
  adj[434] = 1; 
  adj[441] = 1; 
  adj[454] = 1; 
  adj[456] = 1; 
  adj[519] = 1; 
  adj[521] = 1; 
  adj[584] = 1; 
  adj[586] = 1; 
  adj[649] = 1; 
  adj[651] = 1; 
  adj[714] = 1; 
  adj[716] = 1; 
  adj[779] = 1; 
  adj[781] = 1; 
  adj[802] = 1; 
  adj[834] = 1; 
  adj[836] = 1; 
  adj[844] = 1; 
  adj[846] = 1; 
  adj[909] = 1; 
  adj[911] = 1; 
  adj[974] = 1; 
  adj[976] = 1; 
  adj[1027] = 1; 
  adj[1039] = 1; 
  adj[1041] = 1; 
  adj[1104] = 1; 
  adj[1106] = 1; 
  adj[1169] = 1; 
  adj[1171] = 1; 
  adj[1234] = 1; 
  adj[1236] = 1; 
  adj[1261] = 1; 
  adj[1279] = 1; 
  adj[1299] = 1; 
  adj[1301] = 1; 
  adj[1364] = 1; 
  adj[1366] = 1; 
  adj[1404] = 1; 
  adj[1429] = 1; 
  adj[1431] = 1; 
  adj[1494] = 1; 
  adj[1496] = 1; 
  adj[1500] = 1; 
  adj[1559] = 1; 
  adj[1561] = 1; 
  adj[1624] = 1; 
  adj[1626] = 1; 
  adj[1689] = 1; 
  adj[1691] = 1; 
  adj[1754] = 1; 
  adj[1756] = 1; 
  adj[1815] = 1; 
  adj[1819] = 1; 
  adj[1821] = 1; 
  adj[1856] = 1; 
  adj[1884] = 1; 
  adj[1886] = 1; 
  adj[1903] = 1; 
  adj[1949] = 1; 
  adj[1951] = 1; 
  adj[1977] = 1; 
  adj[2014] = 1; 
  adj[2016] = 1; 
  adj[2079] = 1; 
  adj[2081] = 1; 
  adj[2144] = 1; 
  adj[2146] = 1; 
  adj[2188] = 1; 
  adj[2209] = 1; 
  adj[2211] = 1; 
  adj[2274] = 1; 
  adj[2276] = 1; 
  adj[2339] = 1; 
  adj[2341] = 1; 
  adj[2404] = 1; 
  adj[2406] = 1; 
  adj[2469] = 1; 
  adj[2471] = 1; 
  adj[2534] = 1; 
  adj[2536] = 1; 
  adj[2599] = 1; 
  adj[2601] = 1; 
  adj[2664] = 1; 
  adj[2666] = 1; 
  adj[2729] = 1; 
  adj[2731] = 1; 
  adj[2794] = 1; 
  adj[2796] = 1; 
  adj[2821] = 1; 
  adj[2859] = 1; 
  adj[2861] = 1; 
  adj[2899] = 1; 
  adj[2924] = 1; 
  adj[2926] = 1; 
  adj[2989] = 1; 
  adj[2991] = 1; 
  adj[3037] = 1; 
  adj[3054] = 1; 
  adj[3056] = 1; 
  adj[3119] = 1; 
  adj[3121] = 1; 
  adj[3184] = 1; 
  adj[3186] = 1; 
  adj[3206] = 1; 
  adj[3249] = 1; 
  adj[3251] = 1; 
  adj[3314] = 1; 
  adj[3316] = 1; 
  adj[3379] = 1; 
  adj[3381] = 1; 
  adj[3444] = 1; 
  adj[3446] = 1; 
  adj[3509] = 1; 
  adj[3511] = 1; 
  adj[3574] = 1; 
  adj[3576] = 1; 
  adj[3639] = 1; 
  adj[3641] = 1; 
  adj[3647] = 1; 
  adj[3654] = 1; 
  adj[3678] = 1; 
  adj[3704] = 1; 
  adj[3706] = 1; 
  adj[3769] = 1; 
  adj[3771] = 1; 
  adj[3834] = 1; 
  adj[3836] = 1; 
  adj[3861] = 1; 
  adj[3899] = 1; 
  adj[3901] = 1; 
  adj[3964] = 1; 
  adj[3966] = 1; 
  adj[4029] = 1; 
  adj[4031] = 1; 
  adj[4032] = 1; 
  adj[4051] = 1; 
  adj[4088] = 1; 
  adj[4094] = 1; 
  nodeWeight[1*WIDTH-1:0*WIDTH] =  16'h5555; 
  nodeWeight[2*WIDTH-1:1*WIDTH] =  16'h8000; 
  nodeWeight[3*WIDTH-1:2*WIDTH] =  16'h5555; 
  nodeWeight[4*WIDTH-1:3*WIDTH] =  16'h5555; 
  nodeWeight[5*WIDTH-1:4*WIDTH] =  16'h5555; 
  nodeWeight[6*WIDTH-1:5*WIDTH] =  16'h5555; 
  nodeWeight[7*WIDTH-1:6*WIDTH] =  16'h4000; 
  nodeWeight[8*WIDTH-1:7*WIDTH] =  16'h8000; 
  nodeWeight[9*WIDTH-1:8*WIDTH] =  16'h8000; 
  nodeWeight[10*WIDTH-1:9*WIDTH] =  16'h8000; 
  nodeWeight[11*WIDTH-1:10*WIDTH] =  16'h8000; 
  nodeWeight[12*WIDTH-1:11*WIDTH] =  16'h8000; 
  nodeWeight[13*WIDTH-1:12*WIDTH] =  16'h5555; 
  nodeWeight[14*WIDTH-1:13*WIDTH] =  16'h4000; 
  nodeWeight[15*WIDTH-1:14*WIDTH] =  16'h8000; 
  nodeWeight[16*WIDTH-1:15*WIDTH] =  16'h8000; 
  nodeWeight[17*WIDTH-1:16*WIDTH] =  16'h5555; 
  nodeWeight[18*WIDTH-1:17*WIDTH] =  16'h8000; 
  nodeWeight[19*WIDTH-1:18*WIDTH] =  16'h8000; 
  nodeWeight[20*WIDTH-1:19*WIDTH] =  16'h4000; 
  nodeWeight[21*WIDTH-1:20*WIDTH] =  16'h8000; 
  nodeWeight[22*WIDTH-1:21*WIDTH] =  16'h5555; 
  nodeWeight[23*WIDTH-1:22*WIDTH] =  16'h8000; 
  nodeWeight[24*WIDTH-1:23*WIDTH] =  16'h5555; 
  nodeWeight[25*WIDTH-1:24*WIDTH] =  16'h8000; 
  nodeWeight[26*WIDTH-1:25*WIDTH] =  16'h8000; 
  nodeWeight[27*WIDTH-1:26*WIDTH] =  16'h8000; 
  nodeWeight[28*WIDTH-1:27*WIDTH] =  16'h8000; 
  nodeWeight[29*WIDTH-1:28*WIDTH] =  16'h5555; 
  nodeWeight[30*WIDTH-1:29*WIDTH] =  16'h4000; 
  nodeWeight[31*WIDTH-1:30*WIDTH] =  16'h5555; 
  nodeWeight[32*WIDTH-1:31*WIDTH] =  16'h8000; 
  nodeWeight[33*WIDTH-1:32*WIDTH] =  16'h8000; 
  nodeWeight[34*WIDTH-1:33*WIDTH] =  16'h8000; 
  nodeWeight[35*WIDTH-1:34*WIDTH] =  16'h5555; 
  nodeWeight[36*WIDTH-1:35*WIDTH] =  16'h8000; 
  nodeWeight[37*WIDTH-1:36*WIDTH] =  16'h8000; 
  nodeWeight[38*WIDTH-1:37*WIDTH] =  16'h8000; 
  nodeWeight[39*WIDTH-1:38*WIDTH] =  16'h8000; 
  nodeWeight[40*WIDTH-1:39*WIDTH] =  16'h8000; 
  nodeWeight[41*WIDTH-1:40*WIDTH] =  16'h8000; 
  nodeWeight[42*WIDTH-1:41*WIDTH] =  16'h8000; 
  nodeWeight[43*WIDTH-1:42*WIDTH] =  16'h8000; 
  nodeWeight[44*WIDTH-1:43*WIDTH] =  16'h8000; 
  nodeWeight[45*WIDTH-1:44*WIDTH] =  16'h5555; 
  nodeWeight[46*WIDTH-1:45*WIDTH] =  16'h5555; 
  nodeWeight[47*WIDTH-1:46*WIDTH] =  16'h8000; 
  nodeWeight[48*WIDTH-1:47*WIDTH] =  16'h5555; 
  nodeWeight[49*WIDTH-1:48*WIDTH] =  16'h8000; 
  nodeWeight[50*WIDTH-1:49*WIDTH] =  16'h8000; 
  nodeWeight[51*WIDTH-1:50*WIDTH] =  16'h5555; 
  nodeWeight[52*WIDTH-1:51*WIDTH] =  16'h8000; 
  nodeWeight[53*WIDTH-1:52*WIDTH] =  16'h8000; 
  nodeWeight[54*WIDTH-1:53*WIDTH] =  16'h8000; 
  nodeWeight[55*WIDTH-1:54*WIDTH] =  16'h8000; 
  nodeWeight[56*WIDTH-1:55*WIDTH] =  16'h8000; 
  nodeWeight[57*WIDTH-1:56*WIDTH] =  16'h5555; 
  nodeWeight[58*WIDTH-1:57*WIDTH] =  16'h4000; 
  nodeWeight[59*WIDTH-1:58*WIDTH] =  16'h8000; 
  nodeWeight[60*WIDTH-1:59*WIDTH] =  16'h8000; 
  nodeWeight[61*WIDTH-1:60*WIDTH] =  16'h5555; 
  nodeWeight[62*WIDTH-1:61*WIDTH] =  16'h8000; 
  nodeWeight[63*WIDTH-1:62*WIDTH] =  16'h8000; 
  nodeWeight[64*WIDTH-1:63*WIDTH] =  16'h4000; 
  #2 reset = 0;
 end 
 endmodule 
