module pageRank_tb;

localparam N=64;
localparam WIDTH=32;

reg clk;
reg reset;

always begin
  #1 clk  = 1;
  #1 clk = 0;
end

reg [N*N-1:0] adj;
reg [N*WIDTH-1:0] nodeWeight;

reg [5:0] query;
reg [WIDTH+5:0] response;

wire [5:0] request;
wire [WIDTH-1:0] reply;
wire [WIDTH-1:0] node0Val;
// wire [WIDTH-1:0] node1Val;
// wire [WIDTH-1:0] node2Val;
// wire [WIDTH-1:0] node3Val;

// ant  #(N,N,WIDTH) ant(clk,reset,adj,nodeWeight,2'b0,
// 	query,response,
// 	request,reply,node0Val);

//pageRank16 #(N,WIDTH) pr(clk,reset,adj,nodeWeight,node0Val);
//pageRank16V3 #(N,WIDTH) pr(clk,reset,adj,nodeWeight,node0Val);
// pageRankv1 #(N,WIDTH) prv1(clk,reset,adj,nodeWeight,node0Val);
pageRank #(N,WIDTH) prv1(clk,reset,adj,nodeWeight,node0Val);
integer i,j;
initial begin
	reset = 1'b0;

	
	$monitor($time,"node0Val=%d",node0Val);

	#1 reset = 1'b1;


  adj[0] = 0; 
  adj[1] = 1; 
  adj[2] = 0; 
  adj[3] = 0; 
  adj[4] = 0; 
  adj[5] = 0; 
  adj[6] = 0; 
  adj[7] = 0; 
  adj[8] = 0; 
  adj[9] = 0; 
  adj[10] = 0; 
  adj[11] = 0; 
  adj[12] = 0; 
  adj[13] = 0; 
  adj[14] = 0; 
  adj[15] = 0; 
  adj[16] = 0; 
  adj[17] = 0; 
  adj[18] = 0; 
  adj[19] = 0; 
  adj[20] = 0; 
  adj[21] = 0; 
  adj[22] = 0; 
  adj[23] = 0; 
  adj[24] = 0; 
  adj[25] = 0; 
  adj[26] = 0; 
  adj[27] = 0; 
  adj[28] = 0; 
  adj[29] = 0; 
  adj[30] = 0; 
  adj[31] = 0; 
  adj[32] = 0; 
  adj[33] = 0; 
  adj[34] = 0; 
  adj[35] = 0; 
  adj[36] = 0; 
  adj[37] = 0; 
  adj[38] = 0; 
  adj[39] = 0; 
  adj[40] = 0; 
  adj[41] = 0; 
  adj[42] = 0; 
  adj[43] = 0; 
  adj[44] = 0; 
  adj[45] = 0; 
  adj[46] = 0; 
  adj[47] = 0; 
  adj[48] = 0; 
  adj[49] = 0; 
  adj[50] = 0; 
  adj[51] = 0; 
  adj[52] = 0; 
  adj[53] = 0; 
  adj[54] = 0; 
  adj[55] = 0; 
  adj[56] = 0; 
  adj[57] = 0; 
  adj[58] = 0; 
  adj[59] = 0; 
  adj[60] = 0; 
  adj[61] = 0; 
  adj[62] = 0; 
  adj[63] = 1; 
  adj[64] = 1; 
  adj[65] = 0; 
  adj[66] = 1; 
  adj[67] = 0; 
  adj[68] = 0; 
  adj[69] = 0; 
  adj[70] = 0; 
  adj[71] = 0; 
  adj[72] = 0; 
  adj[73] = 0; 
  adj[74] = 0; 
  adj[75] = 0; 
  adj[76] = 0; 
  adj[77] = 0; 
  adj[78] = 0; 
  adj[79] = 0; 
  adj[80] = 0; 
  adj[81] = 0; 
  adj[82] = 0; 
  adj[83] = 0; 
  adj[84] = 0; 
  adj[85] = 0; 
  adj[86] = 0; 
  adj[87] = 0; 
  adj[88] = 0; 
  adj[89] = 0; 
  adj[90] = 0; 
  adj[91] = 0; 
  adj[92] = 0; 
  adj[93] = 0; 
  adj[94] = 0; 
  adj[95] = 0; 
  adj[96] = 0; 
  adj[97] = 0; 
  adj[98] = 0; 
  adj[99] = 0; 
  adj[100] = 0; 
  adj[101] = 0; 
  adj[102] = 0; 
  adj[103] = 0; 
  adj[104] = 0; 
  adj[105] = 0; 
  adj[106] = 0; 
  adj[107] = 0; 
  adj[108] = 0; 
  adj[109] = 0; 
  adj[110] = 0; 
  adj[111] = 0; 
  adj[112] = 0; 
  adj[113] = 0; 
  adj[114] = 0; 
  adj[115] = 0; 
  adj[116] = 0; 
  adj[117] = 0; 
  adj[118] = 0; 
  adj[119] = 0; 
  adj[120] = 0; 
  adj[121] = 0; 
  adj[122] = 0; 
  adj[123] = 0; 
  adj[124] = 0; 
  adj[125] = 0; 
  adj[126] = 0; 
  adj[127] = 0; 
  adj[128] = 0; 
  adj[129] = 1; 
  adj[130] = 0; 
  adj[131] = 1; 
  adj[132] = 0; 
  adj[133] = 0; 
  adj[134] = 0; 
  adj[135] = 0; 
  adj[136] = 0; 
  adj[137] = 0; 
  adj[138] = 0; 
  adj[139] = 0; 
  adj[140] = 0; 
  adj[141] = 0; 
  adj[142] = 0; 
  adj[143] = 0; 
  adj[144] = 0; 
  adj[145] = 0; 
  adj[146] = 0; 
  adj[147] = 0; 
  adj[148] = 0; 
  adj[149] = 0; 
  adj[150] = 0; 
  adj[151] = 0; 
  adj[152] = 0; 
  adj[153] = 0; 
  adj[154] = 0; 
  adj[155] = 0; 
  adj[156] = 0; 
  adj[157] = 0; 
  adj[158] = 0; 
  adj[159] = 0; 
  adj[160] = 0; 
  adj[161] = 0; 
  adj[162] = 0; 
  adj[163] = 0; 
  adj[164] = 0; 
  adj[165] = 0; 
  adj[166] = 0; 
  adj[167] = 0; 
  adj[168] = 0; 
  adj[169] = 0; 
  adj[170] = 0; 
  adj[171] = 0; 
  adj[172] = 0; 
  adj[173] = 0; 
  adj[174] = 0; 
  adj[175] = 0; 
  adj[176] = 0; 
  adj[177] = 0; 
  adj[178] = 0; 
  adj[179] = 0; 
  adj[180] = 0; 
  adj[181] = 0; 
  adj[182] = 0; 
  adj[183] = 0; 
  adj[184] = 0; 
  adj[185] = 0; 
  adj[186] = 0; 
  adj[187] = 0; 
  adj[188] = 0; 
  adj[189] = 0; 
  adj[190] = 0; 
  adj[191] = 0; 
  adj[192] = 0; 
  adj[193] = 0; 
  adj[194] = 1; 
  adj[195] = 0; 
  adj[196] = 1; 
  adj[197] = 0; 
  adj[198] = 0; 
  adj[199] = 0; 
  adj[200] = 0; 
  adj[201] = 0; 
  adj[202] = 0; 
  adj[203] = 0; 
  adj[204] = 0; 
  adj[205] = 0; 
  adj[206] = 0; 
  adj[207] = 0; 
  adj[208] = 0; 
  adj[209] = 0; 
  adj[210] = 0; 
  adj[211] = 0; 
  adj[212] = 0; 
  adj[213] = 0; 
  adj[214] = 0; 
  adj[215] = 0; 
  adj[216] = 0; 
  adj[217] = 0; 
  adj[218] = 0; 
  adj[219] = 0; 
  adj[220] = 0; 
  adj[221] = 0; 
  adj[222] = 0; 
  adj[223] = 0; 
  adj[224] = 0; 
  adj[225] = 0; 
  adj[226] = 0; 
  adj[227] = 0; 
  adj[228] = 0; 
  adj[229] = 0; 
  adj[230] = 0; 
  adj[231] = 0; 
  adj[232] = 0; 
  adj[233] = 0; 
  adj[234] = 0; 
  adj[235] = 0; 
  adj[236] = 0; 
  adj[237] = 0; 
  adj[238] = 0; 
  adj[239] = 0; 
  adj[240] = 0; 
  adj[241] = 0; 
  adj[242] = 0; 
  adj[243] = 0; 
  adj[244] = 0; 
  adj[245] = 0; 
  adj[246] = 0; 
  adj[247] = 0; 
  adj[248] = 0; 
  adj[249] = 0; 
  adj[250] = 0; 
  adj[251] = 0; 
  adj[252] = 0; 
  adj[253] = 0; 
  adj[254] = 0; 
  adj[255] = 0; 
  adj[256] = 0; 
  adj[257] = 0; 
  adj[258] = 0; 
  adj[259] = 1; 
  adj[260] = 0; 
  adj[261] = 1; 
  adj[262] = 0; 
  adj[263] = 0; 
  adj[264] = 0; 
  adj[265] = 0; 
  adj[266] = 0; 
  adj[267] = 0; 
  adj[268] = 0; 
  adj[269] = 0; 
  adj[270] = 0; 
  adj[271] = 0; 
  adj[272] = 0; 
  adj[273] = 0; 
  adj[274] = 0; 
  adj[275] = 0; 
  adj[276] = 0; 
  adj[277] = 0; 
  adj[278] = 0; 
  adj[279] = 0; 
  adj[280] = 0; 
  adj[281] = 0; 
  adj[282] = 0; 
  adj[283] = 0; 
  adj[284] = 0; 
  adj[285] = 0; 
  adj[286] = 0; 
  adj[287] = 0; 
  adj[288] = 0; 
  adj[289] = 0; 
  adj[290] = 0; 
  adj[291] = 0; 
  adj[292] = 0; 
  adj[293] = 0; 
  adj[294] = 0; 
  adj[295] = 0; 
  adj[296] = 0; 
  adj[297] = 0; 
  adj[298] = 0; 
  adj[299] = 0; 
  adj[300] = 0; 
  adj[301] = 0; 
  adj[302] = 0; 
  adj[303] = 0; 
  adj[304] = 0; 
  adj[305] = 0; 
  adj[306] = 0; 
  adj[307] = 0; 
  adj[308] = 0; 
  adj[309] = 0; 
  adj[310] = 0; 
  adj[311] = 0; 
  adj[312] = 0; 
  adj[313] = 0; 
  adj[314] = 0; 
  adj[315] = 0; 
  adj[316] = 0; 
  adj[317] = 0; 
  adj[318] = 0; 
  adj[319] = 0; 
  adj[320] = 0; 
  adj[321] = 0; 
  adj[322] = 0; 
  adj[323] = 0; 
  adj[324] = 1; 
  adj[325] = 0; 
  adj[326] = 1; 
  adj[327] = 0; 
  adj[328] = 0; 
  adj[329] = 0; 
  adj[330] = 0; 
  adj[331] = 0; 
  adj[332] = 0; 
  adj[333] = 0; 
  adj[334] = 0; 
  adj[335] = 0; 
  adj[336] = 0; 
  adj[337] = 0; 
  adj[338] = 0; 
  adj[339] = 0; 
  adj[340] = 0; 
  adj[341] = 0; 
  adj[342] = 0; 
  adj[343] = 0; 
  adj[344] = 0; 
  adj[345] = 0; 
  adj[346] = 0; 
  adj[347] = 0; 
  adj[348] = 0; 
  adj[349] = 0; 
  adj[350] = 0; 
  adj[351] = 0; 
  adj[352] = 0; 
  adj[353] = 0; 
  adj[354] = 0; 
  adj[355] = 0; 
  adj[356] = 0; 
  adj[357] = 0; 
  adj[358] = 0; 
  adj[359] = 0; 
  adj[360] = 0; 
  adj[361] = 0; 
  adj[362] = 0; 
  adj[363] = 0; 
  adj[364] = 0; 
  adj[365] = 0; 
  adj[366] = 0; 
  adj[367] = 0; 
  adj[368] = 0; 
  adj[369] = 0; 
  adj[370] = 0; 
  adj[371] = 0; 
  adj[372] = 0; 
  adj[373] = 0; 
  adj[374] = 0; 
  adj[375] = 0; 
  adj[376] = 0; 
  adj[377] = 0; 
  adj[378] = 0; 
  adj[379] = 0; 
  adj[380] = 0; 
  adj[381] = 0; 
  adj[382] = 0; 
  adj[383] = 0; 
  adj[384] = 0; 
  adj[385] = 0; 
  adj[386] = 0; 
  adj[387] = 0; 
  adj[388] = 0; 
  adj[389] = 1; 
  adj[390] = 0; 
  adj[391] = 1; 
  adj[392] = 0; 
  adj[393] = 0; 
  adj[394] = 0; 
  adj[395] = 0; 
  adj[396] = 0; 
  adj[397] = 0; 
  adj[398] = 0; 
  adj[399] = 0; 
  adj[400] = 0; 
  adj[401] = 0; 
  adj[402] = 0; 
  adj[403] = 0; 
  adj[404] = 0; 
  adj[405] = 0; 
  adj[406] = 0; 
  adj[407] = 0; 
  adj[408] = 0; 
  adj[409] = 0; 
  adj[410] = 0; 
  adj[411] = 0; 
  adj[412] = 0; 
  adj[413] = 0; 
  adj[414] = 0; 
  adj[415] = 0; 
  adj[416] = 0; 
  adj[417] = 0; 
  adj[418] = 0; 
  adj[419] = 0; 
  adj[420] = 0; 
  adj[421] = 0; 
  adj[422] = 0; 
  adj[423] = 0; 
  adj[424] = 0; 
  adj[425] = 0; 
  adj[426] = 0; 
  adj[427] = 0; 
  adj[428] = 0; 
  adj[429] = 0; 
  adj[430] = 0; 
  adj[431] = 0; 
  adj[432] = 0; 
  adj[433] = 0; 
  adj[434] = 0; 
  adj[435] = 0; 
  adj[436] = 0; 
  adj[437] = 0; 
  adj[438] = 0; 
  adj[439] = 0; 
  adj[440] = 0; 
  adj[441] = 0; 
  adj[442] = 0; 
  adj[443] = 0; 
  adj[444] = 0; 
  adj[445] = 0; 
  adj[446] = 0; 
  adj[447] = 0; 
  adj[448] = 0; 
  adj[449] = 0; 
  adj[450] = 0; 
  adj[451] = 0; 
  adj[452] = 0; 
  adj[453] = 0; 
  adj[454] = 1; 
  adj[455] = 0; 
  adj[456] = 1; 
  adj[457] = 0; 
  adj[458] = 0; 
  adj[459] = 0; 
  adj[460] = 0; 
  adj[461] = 0; 
  adj[462] = 0; 
  adj[463] = 0; 
  adj[464] = 0; 
  adj[465] = 0; 
  adj[466] = 0; 
  adj[467] = 0; 
  adj[468] = 0; 
  adj[469] = 0; 
  adj[470] = 0; 
  adj[471] = 0; 
  adj[472] = 0; 
  adj[473] = 0; 
  adj[474] = 0; 
  adj[475] = 0; 
  adj[476] = 0; 
  adj[477] = 0; 
  adj[478] = 0; 
  adj[479] = 0; 
  adj[480] = 0; 
  adj[481] = 0; 
  adj[482] = 0; 
  adj[483] = 0; 
  adj[484] = 0; 
  adj[485] = 0; 
  adj[486] = 0; 
  adj[487] = 0; 
  adj[488] = 0; 
  adj[489] = 0; 
  adj[490] = 0; 
  adj[491] = 0; 
  adj[492] = 0; 
  adj[493] = 0; 
  adj[494] = 0; 
  adj[495] = 0; 
  adj[496] = 0; 
  adj[497] = 0; 
  adj[498] = 0; 
  adj[499] = 0; 
  adj[500] = 0; 
  adj[501] = 0; 
  adj[502] = 0; 
  adj[503] = 0; 
  adj[504] = 0; 
  adj[505] = 0; 
  adj[506] = 0; 
  adj[507] = 0; 
  adj[508] = 0; 
  adj[509] = 0; 
  adj[510] = 0; 
  adj[511] = 0; 
  adj[512] = 0; 
  adj[513] = 0; 
  adj[514] = 0; 
  adj[515] = 0; 
  adj[516] = 0; 
  adj[517] = 0; 
  adj[518] = 0; 
  adj[519] = 1; 
  adj[520] = 0; 
  adj[521] = 1; 
  adj[522] = 0; 
  adj[523] = 0; 
  adj[524] = 0; 
  adj[525] = 0; 
  adj[526] = 0; 
  adj[527] = 0; 
  adj[528] = 0; 
  adj[529] = 0; 
  adj[530] = 0; 
  adj[531] = 0; 
  adj[532] = 0; 
  adj[533] = 0; 
  adj[534] = 0; 
  adj[535] = 0; 
  adj[536] = 0; 
  adj[537] = 0; 
  adj[538] = 0; 
  adj[539] = 0; 
  adj[540] = 0; 
  adj[541] = 0; 
  adj[542] = 0; 
  adj[543] = 0; 
  adj[544] = 0; 
  adj[545] = 0; 
  adj[546] = 0; 
  adj[547] = 0; 
  adj[548] = 0; 
  adj[549] = 0; 
  adj[550] = 0; 
  adj[551] = 0; 
  adj[552] = 0; 
  adj[553] = 0; 
  adj[554] = 0; 
  adj[555] = 0; 
  adj[556] = 0; 
  adj[557] = 0; 
  adj[558] = 0; 
  adj[559] = 0; 
  adj[560] = 0; 
  adj[561] = 0; 
  adj[562] = 0; 
  adj[563] = 0; 
  adj[564] = 0; 
  adj[565] = 0; 
  adj[566] = 0; 
  adj[567] = 0; 
  adj[568] = 0; 
  adj[569] = 0; 
  adj[570] = 0; 
  adj[571] = 0; 
  adj[572] = 0; 
  adj[573] = 0; 
  adj[574] = 0; 
  adj[575] = 0; 
  adj[576] = 0; 
  adj[577] = 0; 
  adj[578] = 0; 
  adj[579] = 0; 
  adj[580] = 0; 
  adj[581] = 0; 
  adj[582] = 0; 
  adj[583] = 0; 
  adj[584] = 1; 
  adj[585] = 0; 
  adj[586] = 1; 
  adj[587] = 0; 
  adj[588] = 0; 
  adj[589] = 0; 
  adj[590] = 0; 
  adj[591] = 0; 
  adj[592] = 0; 
  adj[593] = 0; 
  adj[594] = 0; 
  adj[595] = 0; 
  adj[596] = 0; 
  adj[597] = 0; 
  adj[598] = 0; 
  adj[599] = 0; 
  adj[600] = 0; 
  adj[601] = 0; 
  adj[602] = 0; 
  adj[603] = 0; 
  adj[604] = 0; 
  adj[605] = 0; 
  adj[606] = 0; 
  adj[607] = 0; 
  adj[608] = 0; 
  adj[609] = 0; 
  adj[610] = 0; 
  adj[611] = 0; 
  adj[612] = 0; 
  adj[613] = 0; 
  adj[614] = 0; 
  adj[615] = 0; 
  adj[616] = 0; 
  adj[617] = 0; 
  adj[618] = 0; 
  adj[619] = 0; 
  adj[620] = 0; 
  adj[621] = 0; 
  adj[622] = 0; 
  adj[623] = 0; 
  adj[624] = 0; 
  adj[625] = 0; 
  adj[626] = 0; 
  adj[627] = 0; 
  adj[628] = 0; 
  adj[629] = 0; 
  adj[630] = 0; 
  adj[631] = 0; 
  adj[632] = 0; 
  adj[633] = 0; 
  adj[634] = 0; 
  adj[635] = 0; 
  adj[636] = 0; 
  adj[637] = 0; 
  adj[638] = 0; 
  adj[639] = 0; 
  adj[640] = 0; 
  adj[641] = 0; 
  adj[642] = 0; 
  adj[643] = 0; 
  adj[644] = 0; 
  adj[645] = 0; 
  adj[646] = 0; 
  adj[647] = 0; 
  adj[648] = 0; 
  adj[649] = 1; 
  adj[650] = 0; 
  adj[651] = 1; 
  adj[652] = 0; 
  adj[653] = 0; 
  adj[654] = 0; 
  adj[655] = 0; 
  adj[656] = 0; 
  adj[657] = 0; 
  adj[658] = 0; 
  adj[659] = 0; 
  adj[660] = 0; 
  adj[661] = 0; 
  adj[662] = 0; 
  adj[663] = 0; 
  adj[664] = 0; 
  adj[665] = 0; 
  adj[666] = 0; 
  adj[667] = 0; 
  adj[668] = 0; 
  adj[669] = 0; 
  adj[670] = 0; 
  adj[671] = 0; 
  adj[672] = 0; 
  adj[673] = 0; 
  adj[674] = 0; 
  adj[675] = 0; 
  adj[676] = 0; 
  adj[677] = 0; 
  adj[678] = 0; 
  adj[679] = 0; 
  adj[680] = 0; 
  adj[681] = 0; 
  adj[682] = 0; 
  adj[683] = 0; 
  adj[684] = 0; 
  adj[685] = 0; 
  adj[686] = 0; 
  adj[687] = 0; 
  adj[688] = 0; 
  adj[689] = 0; 
  adj[690] = 0; 
  adj[691] = 0; 
  adj[692] = 0; 
  adj[693] = 0; 
  adj[694] = 0; 
  adj[695] = 0; 
  adj[696] = 0; 
  adj[697] = 0; 
  adj[698] = 0; 
  adj[699] = 0; 
  adj[700] = 0; 
  adj[701] = 0; 
  adj[702] = 0; 
  adj[703] = 0; 
  adj[704] = 0; 
  adj[705] = 0; 
  adj[706] = 0; 
  adj[707] = 0; 
  adj[708] = 0; 
  adj[709] = 0; 
  adj[710] = 0; 
  adj[711] = 0; 
  adj[712] = 0; 
  adj[713] = 0; 
  adj[714] = 1; 
  adj[715] = 0; 
  adj[716] = 1; 
  adj[717] = 0; 
  adj[718] = 0; 
  adj[719] = 0; 
  adj[720] = 0; 
  adj[721] = 0; 
  adj[722] = 0; 
  adj[723] = 0; 
  adj[724] = 0; 
  adj[725] = 0; 
  adj[726] = 0; 
  adj[727] = 0; 
  adj[728] = 0; 
  adj[729] = 0; 
  adj[730] = 0; 
  adj[731] = 0; 
  adj[732] = 0; 
  adj[733] = 0; 
  adj[734] = 0; 
  adj[735] = 0; 
  adj[736] = 0; 
  adj[737] = 0; 
  adj[738] = 0; 
  adj[739] = 0; 
  adj[740] = 0; 
  adj[741] = 0; 
  adj[742] = 0; 
  adj[743] = 0; 
  adj[744] = 0; 
  adj[745] = 0; 
  adj[746] = 0; 
  adj[747] = 0; 
  adj[748] = 0; 
  adj[749] = 0; 
  adj[750] = 0; 
  adj[751] = 0; 
  adj[752] = 0; 
  adj[753] = 0; 
  adj[754] = 0; 
  adj[755] = 0; 
  adj[756] = 0; 
  adj[757] = 0; 
  adj[758] = 0; 
  adj[759] = 0; 
  adj[760] = 0; 
  adj[761] = 0; 
  adj[762] = 0; 
  adj[763] = 0; 
  adj[764] = 0; 
  adj[765] = 0; 
  adj[766] = 0; 
  adj[767] = 0; 
  adj[768] = 0; 
  adj[769] = 0; 
  adj[770] = 0; 
  adj[771] = 0; 
  adj[772] = 0; 
  adj[773] = 0; 
  adj[774] = 0; 
  adj[775] = 0; 
  adj[776] = 0; 
  adj[777] = 0; 
  adj[778] = 0; 
  adj[779] = 1; 
  adj[780] = 0; 
  adj[781] = 1; 
  adj[782] = 0; 
  adj[783] = 0; 
  adj[784] = 0; 
  adj[785] = 0; 
  adj[786] = 0; 
  adj[787] = 0; 
  adj[788] = 0; 
  adj[789] = 0; 
  adj[790] = 0; 
  adj[791] = 0; 
  adj[792] = 0; 
  adj[793] = 0; 
  adj[794] = 0; 
  adj[795] = 0; 
  adj[796] = 0; 
  adj[797] = 0; 
  adj[798] = 0; 
  adj[799] = 0; 
  adj[800] = 0; 
  adj[801] = 0; 
  adj[802] = 0; 
  adj[803] = 0; 
  adj[804] = 0; 
  adj[805] = 0; 
  adj[806] = 0; 
  adj[807] = 0; 
  adj[808] = 0; 
  adj[809] = 0; 
  adj[810] = 0; 
  adj[811] = 0; 
  adj[812] = 0; 
  adj[813] = 0; 
  adj[814] = 0; 
  adj[815] = 0; 
  adj[816] = 0; 
  adj[817] = 0; 
  adj[818] = 0; 
  adj[819] = 0; 
  adj[820] = 0; 
  adj[821] = 0; 
  adj[822] = 0; 
  adj[823] = 0; 
  adj[824] = 0; 
  adj[825] = 0; 
  adj[826] = 0; 
  adj[827] = 0; 
  adj[828] = 0; 
  adj[829] = 0; 
  adj[830] = 0; 
  adj[831] = 1; 
  adj[832] = 0; 
  adj[833] = 0; 
  adj[834] = 0; 
  adj[835] = 0; 
  adj[836] = 0; 
  adj[837] = 0; 
  adj[838] = 0; 
  adj[839] = 0; 
  adj[840] = 0; 
  adj[841] = 0; 
  adj[842] = 0; 
  adj[843] = 0; 
  adj[844] = 1; 
  adj[845] = 0; 
  adj[846] = 1; 
  adj[847] = 0; 
  adj[848] = 0; 
  adj[849] = 0; 
  adj[850] = 0; 
  adj[851] = 0; 
  adj[852] = 0; 
  adj[853] = 0; 
  adj[854] = 0; 
  adj[855] = 0; 
  adj[856] = 0; 
  adj[857] = 0; 
  adj[858] = 0; 
  adj[859] = 0; 
  adj[860] = 0; 
  adj[861] = 0; 
  adj[862] = 0; 
  adj[863] = 0; 
  adj[864] = 0; 
  adj[865] = 0; 
  adj[866] = 0; 
  adj[867] = 0; 
  adj[868] = 0; 
  adj[869] = 0; 
  adj[870] = 0; 
  adj[871] = 0; 
  adj[872] = 0; 
  adj[873] = 0; 
  adj[874] = 0; 
  adj[875] = 0; 
  adj[876] = 0; 
  adj[877] = 0; 
  adj[878] = 0; 
  adj[879] = 0; 
  adj[880] = 0; 
  adj[881] = 0; 
  adj[882] = 0; 
  adj[883] = 0; 
  adj[884] = 0; 
  adj[885] = 0; 
  adj[886] = 0; 
  adj[887] = 0; 
  adj[888] = 0; 
  adj[889] = 0; 
  adj[890] = 0; 
  adj[891] = 0; 
  adj[892] = 0; 
  adj[893] = 0; 
  adj[894] = 0; 
  adj[895] = 0; 
  adj[896] = 0; 
  adj[897] = 0; 
  adj[898] = 0; 
  adj[899] = 0; 
  adj[900] = 0; 
  adj[901] = 0; 
  adj[902] = 0; 
  adj[903] = 0; 
  adj[904] = 0; 
  adj[905] = 0; 
  adj[906] = 0; 
  adj[907] = 0; 
  adj[908] = 0; 
  adj[909] = 1; 
  adj[910] = 0; 
  adj[911] = 1; 
  adj[912] = 0; 
  adj[913] = 0; 
  adj[914] = 0; 
  adj[915] = 0; 
  adj[916] = 0; 
  adj[917] = 0; 
  adj[918] = 0; 
  adj[919] = 0; 
  adj[920] = 0; 
  adj[921] = 0; 
  adj[922] = 0; 
  adj[923] = 0; 
  adj[924] = 0; 
  adj[925] = 0; 
  adj[926] = 0; 
  adj[927] = 0; 
  adj[928] = 0; 
  adj[929] = 0; 
  adj[930] = 0; 
  adj[931] = 0; 
  adj[932] = 0; 
  adj[933] = 0; 
  adj[934] = 0; 
  adj[935] = 0; 
  adj[936] = 0; 
  adj[937] = 0; 
  adj[938] = 0; 
  adj[939] = 0; 
  adj[940] = 0; 
  adj[941] = 0; 
  adj[942] = 0; 
  adj[943] = 0; 
  adj[944] = 0; 
  adj[945] = 0; 
  adj[946] = 0; 
  adj[947] = 0; 
  adj[948] = 0; 
  adj[949] = 0; 
  adj[950] = 0; 
  adj[951] = 0; 
  adj[952] = 0; 
  adj[953] = 0; 
  adj[954] = 0; 
  adj[955] = 0; 
  adj[956] = 0; 
  adj[957] = 0; 
  adj[958] = 0; 
  adj[959] = 0; 
  adj[960] = 0; 
  adj[961] = 0; 
  adj[962] = 0; 
  adj[963] = 0; 
  adj[964] = 0; 
  adj[965] = 0; 
  adj[966] = 0; 
  adj[967] = 0; 
  adj[968] = 0; 
  adj[969] = 0; 
  adj[970] = 0; 
  adj[971] = 0; 
  adj[972] = 0; 
  adj[973] = 0; 
  adj[974] = 1; 
  adj[975] = 0; 
  adj[976] = 1; 
  adj[977] = 0; 
  adj[978] = 0; 
  adj[979] = 0; 
  adj[980] = 0; 
  adj[981] = 0; 
  adj[982] = 0; 
  adj[983] = 0; 
  adj[984] = 0; 
  adj[985] = 0; 
  adj[986] = 0; 
  adj[987] = 0; 
  adj[988] = 0; 
  adj[989] = 0; 
  adj[990] = 0; 
  adj[991] = 0; 
  adj[992] = 0; 
  adj[993] = 0; 
  adj[994] = 0; 
  adj[995] = 0; 
  adj[996] = 0; 
  adj[997] = 0; 
  adj[998] = 0; 
  adj[999] = 0; 
  adj[1000] = 0; 
  adj[1001] = 0; 
  adj[1002] = 0; 
  adj[1003] = 0; 
  adj[1004] = 0; 
  adj[1005] = 0; 
  adj[1006] = 0; 
  adj[1007] = 0; 
  adj[1008] = 0; 
  adj[1009] = 0; 
  adj[1010] = 0; 
  adj[1011] = 0; 
  adj[1012] = 0; 
  adj[1013] = 0; 
  adj[1014] = 0; 
  adj[1015] = 0; 
  adj[1016] = 0; 
  adj[1017] = 0; 
  adj[1018] = 0; 
  adj[1019] = 0; 
  adj[1020] = 0; 
  adj[1021] = 0; 
  adj[1022] = 0; 
  adj[1023] = 0; 
  adj[1024] = 0; 
  adj[1025] = 0; 
  adj[1026] = 0; 
  adj[1027] = 0; 
  adj[1028] = 0; 
  adj[1029] = 0; 
  adj[1030] = 0; 
  adj[1031] = 0; 
  adj[1032] = 0; 
  adj[1033] = 0; 
  adj[1034] = 0; 
  adj[1035] = 0; 
  adj[1036] = 0; 
  adj[1037] = 0; 
  adj[1038] = 0; 
  adj[1039] = 1; 
  adj[1040] = 0; 
  adj[1041] = 1; 
  adj[1042] = 0; 
  adj[1043] = 0; 
  adj[1044] = 0; 
  adj[1045] = 0; 
  adj[1046] = 0; 
  adj[1047] = 0; 
  adj[1048] = 0; 
  adj[1049] = 0; 
  adj[1050] = 0; 
  adj[1051] = 0; 
  adj[1052] = 0; 
  adj[1053] = 0; 
  adj[1054] = 0; 
  adj[1055] = 0; 
  adj[1056] = 0; 
  adj[1057] = 0; 
  adj[1058] = 0; 
  adj[1059] = 0; 
  adj[1060] = 0; 
  adj[1061] = 0; 
  adj[1062] = 0; 
  adj[1063] = 0; 
  adj[1064] = 0; 
  adj[1065] = 0; 
  adj[1066] = 0; 
  adj[1067] = 0; 
  adj[1068] = 0; 
  adj[1069] = 0; 
  adj[1070] = 0; 
  adj[1071] = 0; 
  adj[1072] = 0; 
  adj[1073] = 0; 
  adj[1074] = 0; 
  adj[1075] = 0; 
  adj[1076] = 0; 
  adj[1077] = 0; 
  adj[1078] = 0; 
  adj[1079] = 0; 
  adj[1080] = 0; 
  adj[1081] = 0; 
  adj[1082] = 0; 
  adj[1083] = 0; 
  adj[1084] = 0; 
  adj[1085] = 0; 
  adj[1086] = 0; 
  adj[1087] = 0; 
  adj[1088] = 0; 
  adj[1089] = 0; 
  adj[1090] = 0; 
  adj[1091] = 0; 
  adj[1092] = 0; 
  adj[1093] = 0; 
  adj[1094] = 0; 
  adj[1095] = 0; 
  adj[1096] = 0; 
  adj[1097] = 0; 
  adj[1098] = 0; 
  adj[1099] = 0; 
  adj[1100] = 0; 
  adj[1101] = 0; 
  adj[1102] = 0; 
  adj[1103] = 0; 
  adj[1104] = 1; 
  adj[1105] = 0; 
  adj[1106] = 1; 
  adj[1107] = 0; 
  adj[1108] = 0; 
  adj[1109] = 0; 
  adj[1110] = 0; 
  adj[1111] = 0; 
  adj[1112] = 0; 
  adj[1113] = 0; 
  adj[1114] = 0; 
  adj[1115] = 0; 
  adj[1116] = 0; 
  adj[1117] = 0; 
  adj[1118] = 0; 
  adj[1119] = 0; 
  adj[1120] = 0; 
  adj[1121] = 0; 
  adj[1122] = 0; 
  adj[1123] = 0; 
  adj[1124] = 0; 
  adj[1125] = 0; 
  adj[1126] = 0; 
  adj[1127] = 0; 
  adj[1128] = 0; 
  adj[1129] = 0; 
  adj[1130] = 0; 
  adj[1131] = 0; 
  adj[1132] = 0; 
  adj[1133] = 0; 
  adj[1134] = 0; 
  adj[1135] = 0; 
  adj[1136] = 0; 
  adj[1137] = 0; 
  adj[1138] = 0; 
  adj[1139] = 0; 
  adj[1140] = 1; 
  adj[1141] = 0; 
  adj[1142] = 0; 
  adj[1143] = 0; 
  adj[1144] = 0; 
  adj[1145] = 0; 
  adj[1146] = 0; 
  adj[1147] = 0; 
  adj[1148] = 0; 
  adj[1149] = 0; 
  adj[1150] = 0; 
  adj[1151] = 0; 
  adj[1152] = 0; 
  adj[1153] = 0; 
  adj[1154] = 0; 
  adj[1155] = 0; 
  adj[1156] = 0; 
  adj[1157] = 0; 
  adj[1158] = 0; 
  adj[1159] = 0; 
  adj[1160] = 0; 
  adj[1161] = 0; 
  adj[1162] = 0; 
  adj[1163] = 0; 
  adj[1164] = 0; 
  adj[1165] = 0; 
  adj[1166] = 0; 
  adj[1167] = 0; 
  adj[1168] = 0; 
  adj[1169] = 1; 
  adj[1170] = 0; 
  adj[1171] = 1; 
  adj[1172] = 0; 
  adj[1173] = 0; 
  adj[1174] = 0; 
  adj[1175] = 0; 
  adj[1176] = 0; 
  adj[1177] = 0; 
  adj[1178] = 0; 
  adj[1179] = 0; 
  adj[1180] = 0; 
  adj[1181] = 0; 
  adj[1182] = 0; 
  adj[1183] = 0; 
  adj[1184] = 0; 
  adj[1185] = 0; 
  adj[1186] = 0; 
  adj[1187] = 0; 
  adj[1188] = 0; 
  adj[1189] = 0; 
  adj[1190] = 0; 
  adj[1191] = 0; 
  adj[1192] = 0; 
  adj[1193] = 0; 
  adj[1194] = 0; 
  adj[1195] = 0; 
  adj[1196] = 0; 
  adj[1197] = 0; 
  adj[1198] = 0; 
  adj[1199] = 0; 
  adj[1200] = 0; 
  adj[1201] = 0; 
  adj[1202] = 0; 
  adj[1203] = 0; 
  adj[1204] = 0; 
  adj[1205] = 0; 
  adj[1206] = 0; 
  adj[1207] = 0; 
  adj[1208] = 0; 
  adj[1209] = 0; 
  adj[1210] = 0; 
  adj[1211] = 0; 
  adj[1212] = 0; 
  adj[1213] = 0; 
  adj[1214] = 0; 
  adj[1215] = 0; 
  adj[1216] = 0; 
  adj[1217] = 0; 
  adj[1218] = 0; 
  adj[1219] = 0; 
  adj[1220] = 0; 
  adj[1221] = 0; 
  adj[1222] = 0; 
  adj[1223] = 0; 
  adj[1224] = 0; 
  adj[1225] = 0; 
  adj[1226] = 0; 
  adj[1227] = 0; 
  adj[1228] = 0; 
  adj[1229] = 0; 
  adj[1230] = 0; 
  adj[1231] = 0; 
  adj[1232] = 0; 
  adj[1233] = 0; 
  adj[1234] = 1; 
  adj[1235] = 0; 
  adj[1236] = 1; 
  adj[1237] = 0; 
  adj[1238] = 0; 
  adj[1239] = 0; 
  adj[1240] = 0; 
  adj[1241] = 0; 
  adj[1242] = 0; 
  adj[1243] = 0; 
  adj[1244] = 0; 
  adj[1245] = 0; 
  adj[1246] = 0; 
  adj[1247] = 0; 
  adj[1248] = 0; 
  adj[1249] = 0; 
  adj[1250] = 0; 
  adj[1251] = 0; 
  adj[1252] = 0; 
  adj[1253] = 0; 
  adj[1254] = 0; 
  adj[1255] = 0; 
  adj[1256] = 0; 
  adj[1257] = 0; 
  adj[1258] = 0; 
  adj[1259] = 0; 
  adj[1260] = 0; 
  adj[1261] = 0; 
  adj[1262] = 0; 
  adj[1263] = 0; 
  adj[1264] = 0; 
  adj[1265] = 0; 
  adj[1266] = 0; 
  adj[1267] = 0; 
  adj[1268] = 0; 
  adj[1269] = 0; 
  adj[1270] = 0; 
  adj[1271] = 0; 
  adj[1272] = 0; 
  adj[1273] = 0; 
  adj[1274] = 0; 
  adj[1275] = 0; 
  adj[1276] = 0; 
  adj[1277] = 0; 
  adj[1278] = 0; 
  adj[1279] = 0; 
  adj[1280] = 0; 
  adj[1281] = 0; 
  adj[1282] = 0; 
  adj[1283] = 0; 
  adj[1284] = 0; 
  adj[1285] = 0; 
  adj[1286] = 0; 
  adj[1287] = 0; 
  adj[1288] = 0; 
  adj[1289] = 0; 
  adj[1290] = 0; 
  adj[1291] = 0; 
  adj[1292] = 0; 
  adj[1293] = 0; 
  adj[1294] = 0; 
  adj[1295] = 0; 
  adj[1296] = 0; 
  adj[1297] = 0; 
  adj[1298] = 0; 
  adj[1299] = 1; 
  adj[1300] = 0; 
  adj[1301] = 1; 
  adj[1302] = 0; 
  adj[1303] = 0; 
  adj[1304] = 0; 
  adj[1305] = 0; 
  adj[1306] = 0; 
  adj[1307] = 0; 
  adj[1308] = 0; 
  adj[1309] = 0; 
  adj[1310] = 0; 
  adj[1311] = 0; 
  adj[1312] = 0; 
  adj[1313] = 0; 
  adj[1314] = 0; 
  adj[1315] = 0; 
  adj[1316] = 0; 
  adj[1317] = 0; 
  adj[1318] = 0; 
  adj[1319] = 0; 
  adj[1320] = 0; 
  adj[1321] = 0; 
  adj[1322] = 0; 
  adj[1323] = 0; 
  adj[1324] = 0; 
  adj[1325] = 0; 
  adj[1326] = 0; 
  adj[1327] = 0; 
  adj[1328] = 0; 
  adj[1329] = 0; 
  adj[1330] = 0; 
  adj[1331] = 0; 
  adj[1332] = 0; 
  adj[1333] = 0; 
  adj[1334] = 0; 
  adj[1335] = 0; 
  adj[1336] = 0; 
  adj[1337] = 0; 
  adj[1338] = 0; 
  adj[1339] = 0; 
  adj[1340] = 0; 
  adj[1341] = 0; 
  adj[1342] = 0; 
  adj[1343] = 0; 
  adj[1344] = 0; 
  adj[1345] = 0; 
  adj[1346] = 0; 
  adj[1347] = 0; 
  adj[1348] = 0; 
  adj[1349] = 0; 
  adj[1350] = 0; 
  adj[1351] = 0; 
  adj[1352] = 0; 
  adj[1353] = 0; 
  adj[1354] = 0; 
  adj[1355] = 0; 
  adj[1356] = 0; 
  adj[1357] = 0; 
  adj[1358] = 0; 
  adj[1359] = 0; 
  adj[1360] = 0; 
  adj[1361] = 0; 
  adj[1362] = 0; 
  adj[1363] = 0; 
  adj[1364] = 1; 
  adj[1365] = 0; 
  adj[1366] = 1; 
  adj[1367] = 0; 
  adj[1368] = 0; 
  adj[1369] = 0; 
  adj[1370] = 0; 
  adj[1371] = 1; 
  adj[1372] = 0; 
  adj[1373] = 0; 
  adj[1374] = 0; 
  adj[1375] = 0; 
  adj[1376] = 0; 
  adj[1377] = 0; 
  adj[1378] = 0; 
  adj[1379] = 0; 
  adj[1380] = 0; 
  adj[1381] = 0; 
  adj[1382] = 0; 
  adj[1383] = 0; 
  adj[1384] = 0; 
  adj[1385] = 0; 
  adj[1386] = 0; 
  adj[1387] = 0; 
  adj[1388] = 0; 
  adj[1389] = 0; 
  adj[1390] = 0; 
  adj[1391] = 0; 
  adj[1392] = 0; 
  adj[1393] = 0; 
  adj[1394] = 0; 
  adj[1395] = 0; 
  adj[1396] = 0; 
  adj[1397] = 0; 
  adj[1398] = 0; 
  adj[1399] = 0; 
  adj[1400] = 0; 
  adj[1401] = 0; 
  adj[1402] = 0; 
  adj[1403] = 0; 
  adj[1404] = 0; 
  adj[1405] = 0; 
  adj[1406] = 0; 
  adj[1407] = 0; 
  adj[1408] = 0; 
  adj[1409] = 0; 
  adj[1410] = 0; 
  adj[1411] = 0; 
  adj[1412] = 0; 
  adj[1413] = 0; 
  adj[1414] = 0; 
  adj[1415] = 0; 
  adj[1416] = 0; 
  adj[1417] = 0; 
  adj[1418] = 0; 
  adj[1419] = 0; 
  adj[1420] = 0; 
  adj[1421] = 0; 
  adj[1422] = 0; 
  adj[1423] = 0; 
  adj[1424] = 0; 
  adj[1425] = 0; 
  adj[1426] = 0; 
  adj[1427] = 0; 
  adj[1428] = 0; 
  adj[1429] = 1; 
  adj[1430] = 0; 
  adj[1431] = 1; 
  adj[1432] = 0; 
  adj[1433] = 0; 
  adj[1434] = 0; 
  adj[1435] = 0; 
  adj[1436] = 0; 
  adj[1437] = 0; 
  adj[1438] = 0; 
  adj[1439] = 0; 
  adj[1440] = 0; 
  adj[1441] = 0; 
  adj[1442] = 0; 
  adj[1443] = 0; 
  adj[1444] = 0; 
  adj[1445] = 0; 
  adj[1446] = 0; 
  adj[1447] = 0; 
  adj[1448] = 0; 
  adj[1449] = 0; 
  adj[1450] = 0; 
  adj[1451] = 0; 
  adj[1452] = 0; 
  adj[1453] = 0; 
  adj[1454] = 0; 
  adj[1455] = 0; 
  adj[1456] = 0; 
  adj[1457] = 0; 
  adj[1458] = 0; 
  adj[1459] = 0; 
  adj[1460] = 0; 
  adj[1461] = 0; 
  adj[1462] = 0; 
  adj[1463] = 0; 
  adj[1464] = 0; 
  adj[1465] = 0; 
  adj[1466] = 0; 
  adj[1467] = 0; 
  adj[1468] = 0; 
  adj[1469] = 0; 
  adj[1470] = 0; 
  adj[1471] = 0; 
  adj[1472] = 0; 
  adj[1473] = 0; 
  adj[1474] = 0; 
  adj[1475] = 0; 
  adj[1476] = 0; 
  adj[1477] = 0; 
  adj[1478] = 0; 
  adj[1479] = 0; 
  adj[1480] = 0; 
  adj[1481] = 0; 
  adj[1482] = 0; 
  adj[1483] = 0; 
  adj[1484] = 0; 
  adj[1485] = 0; 
  adj[1486] = 0; 
  adj[1487] = 0; 
  adj[1488] = 0; 
  adj[1489] = 0; 
  adj[1490] = 0; 
  adj[1491] = 0; 
  adj[1492] = 0; 
  adj[1493] = 0; 
  adj[1494] = 1; 
  adj[1495] = 0; 
  adj[1496] = 1; 
  adj[1497] = 0; 
  adj[1498] = 0; 
  adj[1499] = 0; 
  adj[1500] = 0; 
  adj[1501] = 0; 
  adj[1502] = 0; 
  adj[1503] = 0; 
  adj[1504] = 0; 
  adj[1505] = 0; 
  adj[1506] = 0; 
  adj[1507] = 0; 
  adj[1508] = 0; 
  adj[1509] = 0; 
  adj[1510] = 0; 
  adj[1511] = 0; 
  adj[1512] = 0; 
  adj[1513] = 0; 
  adj[1514] = 0; 
  adj[1515] = 0; 
  adj[1516] = 0; 
  adj[1517] = 0; 
  adj[1518] = 0; 
  adj[1519] = 0; 
  adj[1520] = 0; 
  adj[1521] = 0; 
  adj[1522] = 0; 
  adj[1523] = 0; 
  adj[1524] = 0; 
  adj[1525] = 0; 
  adj[1526] = 0; 
  adj[1527] = 0; 
  adj[1528] = 0; 
  adj[1529] = 0; 
  adj[1530] = 0; 
  adj[1531] = 0; 
  adj[1532] = 0; 
  adj[1533] = 0; 
  adj[1534] = 0; 
  adj[1535] = 0; 
  adj[1536] = 0; 
  adj[1537] = 0; 
  adj[1538] = 0; 
  adj[1539] = 0; 
  adj[1540] = 0; 
  adj[1541] = 0; 
  adj[1542] = 0; 
  adj[1543] = 0; 
  adj[1544] = 0; 
  adj[1545] = 0; 
  adj[1546] = 0; 
  adj[1547] = 0; 
  adj[1548] = 0; 
  adj[1549] = 0; 
  adj[1550] = 0; 
  adj[1551] = 0; 
  adj[1552] = 0; 
  adj[1553] = 0; 
  adj[1554] = 0; 
  adj[1555] = 0; 
  adj[1556] = 0; 
  adj[1557] = 0; 
  adj[1558] = 0; 
  adj[1559] = 1; 
  adj[1560] = 0; 
  adj[1561] = 1; 
  adj[1562] = 0; 
  adj[1563] = 0; 
  adj[1564] = 0; 
  adj[1565] = 0; 
  adj[1566] = 0; 
  adj[1567] = 0; 
  adj[1568] = 0; 
  adj[1569] = 0; 
  adj[1570] = 0; 
  adj[1571] = 0; 
  adj[1572] = 0; 
  adj[1573] = 0; 
  adj[1574] = 0; 
  adj[1575] = 0; 
  adj[1576] = 0; 
  adj[1577] = 0; 
  adj[1578] = 0; 
  adj[1579] = 0; 
  adj[1580] = 0; 
  adj[1581] = 0; 
  adj[1582] = 0; 
  adj[1583] = 0; 
  adj[1584] = 0; 
  adj[1585] = 0; 
  adj[1586] = 0; 
  adj[1587] = 0; 
  adj[1588] = 0; 
  adj[1589] = 0; 
  adj[1590] = 0; 
  adj[1591] = 0; 
  adj[1592] = 0; 
  adj[1593] = 0; 
  adj[1594] = 0; 
  adj[1595] = 0; 
  adj[1596] = 0; 
  adj[1597] = 0; 
  adj[1598] = 0; 
  adj[1599] = 0; 
  adj[1600] = 0; 
  adj[1601] = 0; 
  adj[1602] = 0; 
  adj[1603] = 0; 
  adj[1604] = 0; 
  adj[1605] = 0; 
  adj[1606] = 0; 
  adj[1607] = 0; 
  adj[1608] = 0; 
  adj[1609] = 0; 
  adj[1610] = 0; 
  adj[1611] = 0; 
  adj[1612] = 0; 
  adj[1613] = 0; 
  adj[1614] = 0; 
  adj[1615] = 0; 
  adj[1616] = 0; 
  adj[1617] = 0; 
  adj[1618] = 0; 
  adj[1619] = 0; 
  adj[1620] = 0; 
  adj[1621] = 0; 
  adj[1622] = 0; 
  adj[1623] = 0; 
  adj[1624] = 1; 
  adj[1625] = 0; 
  adj[1626] = 1; 
  adj[1627] = 0; 
  adj[1628] = 0; 
  adj[1629] = 0; 
  adj[1630] = 0; 
  adj[1631] = 0; 
  adj[1632] = 0; 
  adj[1633] = 0; 
  adj[1634] = 0; 
  adj[1635] = 0; 
  adj[1636] = 0; 
  adj[1637] = 0; 
  adj[1638] = 0; 
  adj[1639] = 0; 
  adj[1640] = 0; 
  adj[1641] = 0; 
  adj[1642] = 0; 
  adj[1643] = 0; 
  adj[1644] = 0; 
  adj[1645] = 0; 
  adj[1646] = 0; 
  adj[1647] = 0; 
  adj[1648] = 0; 
  adj[1649] = 0; 
  adj[1650] = 0; 
  adj[1651] = 0; 
  adj[1652] = 0; 
  adj[1653] = 0; 
  adj[1654] = 0; 
  adj[1655] = 0; 
  adj[1656] = 0; 
  adj[1657] = 0; 
  adj[1658] = 0; 
  adj[1659] = 0; 
  adj[1660] = 0; 
  adj[1661] = 0; 
  adj[1662] = 0; 
  adj[1663] = 0; 
  adj[1664] = 0; 
  adj[1665] = 0; 
  adj[1666] = 0; 
  adj[1667] = 0; 
  adj[1668] = 0; 
  adj[1669] = 0; 
  adj[1670] = 0; 
  adj[1671] = 0; 
  adj[1672] = 0; 
  adj[1673] = 0; 
  adj[1674] = 0; 
  adj[1675] = 0; 
  adj[1676] = 0; 
  adj[1677] = 0; 
  adj[1678] = 0; 
  adj[1679] = 0; 
  adj[1680] = 0; 
  adj[1681] = 0; 
  adj[1682] = 0; 
  adj[1683] = 0; 
  adj[1684] = 0; 
  adj[1685] = 0; 
  adj[1686] = 0; 
  adj[1687] = 0; 
  adj[1688] = 0; 
  adj[1689] = 1; 
  adj[1690] = 0; 
  adj[1691] = 1; 
  adj[1692] = 0; 
  adj[1693] = 0; 
  adj[1694] = 0; 
  adj[1695] = 0; 
  adj[1696] = 0; 
  adj[1697] = 0; 
  adj[1698] = 0; 
  adj[1699] = 0; 
  adj[1700] = 0; 
  adj[1701] = 0; 
  adj[1702] = 0; 
  adj[1703] = 0; 
  adj[1704] = 0; 
  adj[1705] = 0; 
  adj[1706] = 0; 
  adj[1707] = 0; 
  adj[1708] = 0; 
  adj[1709] = 0; 
  adj[1710] = 0; 
  adj[1711] = 0; 
  adj[1712] = 0; 
  adj[1713] = 0; 
  adj[1714] = 0; 
  adj[1715] = 0; 
  adj[1716] = 0; 
  adj[1717] = 0; 
  adj[1718] = 0; 
  adj[1719] = 0; 
  adj[1720] = 0; 
  adj[1721] = 0; 
  adj[1722] = 0; 
  adj[1723] = 0; 
  adj[1724] = 0; 
  adj[1725] = 0; 
  adj[1726] = 0; 
  adj[1727] = 0; 
  adj[1728] = 0; 
  adj[1729] = 0; 
  adj[1730] = 0; 
  adj[1731] = 0; 
  adj[1732] = 0; 
  adj[1733] = 0; 
  adj[1734] = 0; 
  adj[1735] = 0; 
  adj[1736] = 0; 
  adj[1737] = 0; 
  adj[1738] = 0; 
  adj[1739] = 0; 
  adj[1740] = 0; 
  adj[1741] = 0; 
  adj[1742] = 0; 
  adj[1743] = 0; 
  adj[1744] = 0; 
  adj[1745] = 0; 
  adj[1746] = 0; 
  adj[1747] = 0; 
  adj[1748] = 0; 
  adj[1749] = 1; 
  adj[1750] = 0; 
  adj[1751] = 0; 
  adj[1752] = 0; 
  adj[1753] = 0; 
  adj[1754] = 1; 
  adj[1755] = 0; 
  adj[1756] = 1; 
  adj[1757] = 0; 
  adj[1758] = 0; 
  adj[1759] = 0; 
  adj[1760] = 0; 
  adj[1761] = 0; 
  adj[1762] = 0; 
  adj[1763] = 0; 
  adj[1764] = 0; 
  adj[1765] = 0; 
  adj[1766] = 0; 
  adj[1767] = 1; 
  adj[1768] = 0; 
  adj[1769] = 0; 
  adj[1770] = 0; 
  adj[1771] = 0; 
  adj[1772] = 0; 
  adj[1773] = 0; 
  adj[1774] = 0; 
  adj[1775] = 0; 
  adj[1776] = 0; 
  adj[1777] = 0; 
  adj[1778] = 0; 
  adj[1779] = 0; 
  adj[1780] = 0; 
  adj[1781] = 0; 
  adj[1782] = 0; 
  adj[1783] = 0; 
  adj[1784] = 0; 
  adj[1785] = 0; 
  adj[1786] = 0; 
  adj[1787] = 0; 
  adj[1788] = 0; 
  adj[1789] = 0; 
  adj[1790] = 0; 
  adj[1791] = 0; 
  adj[1792] = 0; 
  adj[1793] = 0; 
  adj[1794] = 0; 
  adj[1795] = 0; 
  adj[1796] = 0; 
  adj[1797] = 0; 
  adj[1798] = 0; 
  adj[1799] = 0; 
  adj[1800] = 0; 
  adj[1801] = 0; 
  adj[1802] = 0; 
  adj[1803] = 0; 
  adj[1804] = 0; 
  adj[1805] = 0; 
  adj[1806] = 0; 
  adj[1807] = 0; 
  adj[1808] = 0; 
  adj[1809] = 0; 
  adj[1810] = 0; 
  adj[1811] = 0; 
  adj[1812] = 0; 
  adj[1813] = 0; 
  adj[1814] = 0; 
  adj[1815] = 0; 
  adj[1816] = 0; 
  adj[1817] = 0; 
  adj[1818] = 0; 
  adj[1819] = 1; 
  adj[1820] = 0; 
  adj[1821] = 1; 
  adj[1822] = 0; 
  adj[1823] = 0; 
  adj[1824] = 0; 
  adj[1825] = 0; 
  adj[1826] = 0; 
  adj[1827] = 0; 
  adj[1828] = 0; 
  adj[1829] = 0; 
  adj[1830] = 0; 
  adj[1831] = 0; 
  adj[1832] = 0; 
  adj[1833] = 0; 
  adj[1834] = 0; 
  adj[1835] = 0; 
  adj[1836] = 0; 
  adj[1837] = 0; 
  adj[1838] = 0; 
  adj[1839] = 0; 
  adj[1840] = 0; 
  adj[1841] = 0; 
  adj[1842] = 0; 
  adj[1843] = 0; 
  adj[1844] = 0; 
  adj[1845] = 0; 
  adj[1846] = 0; 
  adj[1847] = 0; 
  adj[1848] = 0; 
  adj[1849] = 0; 
  adj[1850] = 0; 
  adj[1851] = 0; 
  adj[1852] = 0; 
  adj[1853] = 0; 
  adj[1854] = 0; 
  adj[1855] = 0; 
  adj[1856] = 0; 
  adj[1857] = 0; 
  adj[1858] = 0; 
  adj[1859] = 0; 
  adj[1860] = 0; 
  adj[1861] = 0; 
  adj[1862] = 0; 
  adj[1863] = 0; 
  adj[1864] = 0; 
  adj[1865] = 0; 
  adj[1866] = 0; 
  adj[1867] = 0; 
  adj[1868] = 0; 
  adj[1869] = 0; 
  adj[1870] = 0; 
  adj[1871] = 0; 
  adj[1872] = 0; 
  adj[1873] = 0; 
  adj[1874] = 0; 
  adj[1875] = 0; 
  adj[1876] = 0; 
  adj[1877] = 0; 
  adj[1878] = 0; 
  adj[1879] = 0; 
  adj[1880] = 0; 
  adj[1881] = 0; 
  adj[1882] = 0; 
  adj[1883] = 0; 
  adj[1884] = 1; 
  adj[1885] = 0; 
  adj[1886] = 1; 
  adj[1887] = 0; 
  adj[1888] = 0; 
  adj[1889] = 0; 
  adj[1890] = 0; 
  adj[1891] = 0; 
  adj[1892] = 0; 
  adj[1893] = 0; 
  adj[1894] = 0; 
  adj[1895] = 0; 
  adj[1896] = 0; 
  adj[1897] = 0; 
  adj[1898] = 0; 
  adj[1899] = 0; 
  adj[1900] = 0; 
  adj[1901] = 0; 
  adj[1902] = 0; 
  adj[1903] = 0; 
  adj[1904] = 0; 
  adj[1905] = 0; 
  adj[1906] = 0; 
  adj[1907] = 0; 
  adj[1908] = 0; 
  adj[1909] = 0; 
  adj[1910] = 0; 
  adj[1911] = 0; 
  adj[1912] = 0; 
  adj[1913] = 0; 
  adj[1914] = 0; 
  adj[1915] = 0; 
  adj[1916] = 0; 
  adj[1917] = 0; 
  adj[1918] = 0; 
  adj[1919] = 0; 
  adj[1920] = 0; 
  adj[1921] = 0; 
  adj[1922] = 0; 
  adj[1923] = 0; 
  adj[1924] = 0; 
  adj[1925] = 0; 
  adj[1926] = 0; 
  adj[1927] = 0; 
  adj[1928] = 0; 
  adj[1929] = 0; 
  adj[1930] = 0; 
  adj[1931] = 0; 
  adj[1932] = 0; 
  adj[1933] = 0; 
  adj[1934] = 0; 
  adj[1935] = 0; 
  adj[1936] = 0; 
  adj[1937] = 0; 
  adj[1938] = 0; 
  adj[1939] = 0; 
  adj[1940] = 0; 
  adj[1941] = 0; 
  adj[1942] = 0; 
  adj[1943] = 0; 
  adj[1944] = 0; 
  adj[1945] = 0; 
  adj[1946] = 0; 
  adj[1947] = 0; 
  adj[1948] = 0; 
  adj[1949] = 1; 
  adj[1950] = 0; 
  adj[1951] = 1; 
  adj[1952] = 0; 
  adj[1953] = 0; 
  adj[1954] = 0; 
  adj[1955] = 0; 
  adj[1956] = 0; 
  adj[1957] = 0; 
  adj[1958] = 0; 
  adj[1959] = 0; 
  adj[1960] = 0; 
  adj[1961] = 0; 
  adj[1962] = 0; 
  adj[1963] = 0; 
  adj[1964] = 0; 
  adj[1965] = 0; 
  adj[1966] = 0; 
  adj[1967] = 0; 
  adj[1968] = 0; 
  adj[1969] = 0; 
  adj[1970] = 0; 
  adj[1971] = 0; 
  adj[1972] = 0; 
  adj[1973] = 0; 
  adj[1974] = 0; 
  adj[1975] = 0; 
  adj[1976] = 0; 
  adj[1977] = 0; 
  adj[1978] = 0; 
  adj[1979] = 0; 
  adj[1980] = 0; 
  adj[1981] = 0; 
  adj[1982] = 0; 
  adj[1983] = 0; 
  adj[1984] = 0; 
  adj[1985] = 0; 
  adj[1986] = 0; 
  adj[1987] = 0; 
  adj[1988] = 0; 
  adj[1989] = 0; 
  adj[1990] = 0; 
  adj[1991] = 0; 
  adj[1992] = 0; 
  adj[1993] = 0; 
  adj[1994] = 0; 
  adj[1995] = 0; 
  adj[1996] = 0; 
  adj[1997] = 0; 
  adj[1998] = 0; 
  adj[1999] = 0; 
  adj[2000] = 0; 
  adj[2001] = 0; 
  adj[2002] = 0; 
  adj[2003] = 0; 
  adj[2004] = 0; 
  adj[2005] = 0; 
  adj[2006] = 0; 
  adj[2007] = 0; 
  adj[2008] = 0; 
  adj[2009] = 0; 
  adj[2010] = 0; 
  adj[2011] = 0; 
  adj[2012] = 0; 
  adj[2013] = 0; 
  adj[2014] = 1; 
  adj[2015] = 0; 
  adj[2016] = 1; 
  adj[2017] = 0; 
  adj[2018] = 0; 
  adj[2019] = 0; 
  adj[2020] = 0; 
  adj[2021] = 0; 
  adj[2022] = 0; 
  adj[2023] = 0; 
  adj[2024] = 0; 
  adj[2025] = 0; 
  adj[2026] = 0; 
  adj[2027] = 0; 
  adj[2028] = 0; 
  adj[2029] = 0; 
  adj[2030] = 0; 
  adj[2031] = 0; 
  adj[2032] = 0; 
  adj[2033] = 0; 
  adj[2034] = 0; 
  adj[2035] = 0; 
  adj[2036] = 0; 
  adj[2037] = 0; 
  adj[2038] = 0; 
  adj[2039] = 0; 
  adj[2040] = 0; 
  adj[2041] = 0; 
  adj[2042] = 0; 
  adj[2043] = 0; 
  adj[2044] = 0; 
  adj[2045] = 0; 
  adj[2046] = 0; 
  adj[2047] = 0; 
  adj[2048] = 0; 
  adj[2049] = 0; 
  adj[2050] = 0; 
  adj[2051] = 0; 
  adj[2052] = 0; 
  adj[2053] = 0; 
  adj[2054] = 0; 
  adj[2055] = 0; 
  adj[2056] = 0; 
  adj[2057] = 0; 
  adj[2058] = 0; 
  adj[2059] = 0; 
  adj[2060] = 0; 
  adj[2061] = 0; 
  adj[2062] = 0; 
  adj[2063] = 0; 
  adj[2064] = 0; 
  adj[2065] = 0; 
  adj[2066] = 0; 
  adj[2067] = 0; 
  adj[2068] = 0; 
  adj[2069] = 0; 
  adj[2070] = 0; 
  adj[2071] = 0; 
  adj[2072] = 0; 
  adj[2073] = 0; 
  adj[2074] = 0; 
  adj[2075] = 0; 
  adj[2076] = 0; 
  adj[2077] = 0; 
  adj[2078] = 0; 
  adj[2079] = 1; 
  adj[2080] = 0; 
  adj[2081] = 1; 
  adj[2082] = 0; 
  adj[2083] = 0; 
  adj[2084] = 0; 
  adj[2085] = 0; 
  adj[2086] = 0; 
  adj[2087] = 0; 
  adj[2088] = 0; 
  adj[2089] = 0; 
  adj[2090] = 0; 
  adj[2091] = 0; 
  adj[2092] = 0; 
  adj[2093] = 0; 
  adj[2094] = 0; 
  adj[2095] = 0; 
  adj[2096] = 0; 
  adj[2097] = 0; 
  adj[2098] = 0; 
  adj[2099] = 0; 
  adj[2100] = 0; 
  adj[2101] = 0; 
  adj[2102] = 0; 
  adj[2103] = 0; 
  adj[2104] = 0; 
  adj[2105] = 0; 
  adj[2106] = 0; 
  adj[2107] = 0; 
  adj[2108] = 0; 
  adj[2109] = 0; 
  adj[2110] = 0; 
  adj[2111] = 0; 
  adj[2112] = 0; 
  adj[2113] = 0; 
  adj[2114] = 0; 
  adj[2115] = 0; 
  adj[2116] = 0; 
  adj[2117] = 0; 
  adj[2118] = 0; 
  adj[2119] = 0; 
  adj[2120] = 0; 
  adj[2121] = 0; 
  adj[2122] = 0; 
  adj[2123] = 0; 
  adj[2124] = 0; 
  adj[2125] = 0; 
  adj[2126] = 0; 
  adj[2127] = 0; 
  adj[2128] = 0; 
  adj[2129] = 0; 
  adj[2130] = 0; 
  adj[2131] = 0; 
  adj[2132] = 0; 
  adj[2133] = 0; 
  adj[2134] = 0; 
  adj[2135] = 0; 
  adj[2136] = 0; 
  adj[2137] = 0; 
  adj[2138] = 0; 
  adj[2139] = 0; 
  adj[2140] = 0; 
  adj[2141] = 0; 
  adj[2142] = 0; 
  adj[2143] = 0; 
  adj[2144] = 1; 
  adj[2145] = 0; 
  adj[2146] = 1; 
  adj[2147] = 0; 
  adj[2148] = 0; 
  adj[2149] = 0; 
  adj[2150] = 0; 
  adj[2151] = 0; 
  adj[2152] = 0; 
  adj[2153] = 0; 
  adj[2154] = 0; 
  adj[2155] = 0; 
  adj[2156] = 0; 
  adj[2157] = 0; 
  adj[2158] = 0; 
  adj[2159] = 0; 
  adj[2160] = 0; 
  adj[2161] = 0; 
  adj[2162] = 0; 
  adj[2163] = 0; 
  adj[2164] = 0; 
  adj[2165] = 0; 
  adj[2166] = 0; 
  adj[2167] = 0; 
  adj[2168] = 0; 
  adj[2169] = 0; 
  adj[2170] = 0; 
  adj[2171] = 0; 
  adj[2172] = 0; 
  adj[2173] = 0; 
  adj[2174] = 0; 
  adj[2175] = 0; 
  adj[2176] = 0; 
  adj[2177] = 0; 
  adj[2178] = 0; 
  adj[2179] = 0; 
  adj[2180] = 0; 
  adj[2181] = 0; 
  adj[2182] = 0; 
  adj[2183] = 0; 
  adj[2184] = 0; 
  adj[2185] = 0; 
  adj[2186] = 0; 
  adj[2187] = 0; 
  adj[2188] = 0; 
  adj[2189] = 0; 
  adj[2190] = 0; 
  adj[2191] = 0; 
  adj[2192] = 0; 
  adj[2193] = 0; 
  adj[2194] = 0; 
  adj[2195] = 0; 
  adj[2196] = 0; 
  adj[2197] = 0; 
  adj[2198] = 0; 
  adj[2199] = 0; 
  adj[2200] = 0; 
  adj[2201] = 0; 
  adj[2202] = 0; 
  adj[2203] = 0; 
  adj[2204] = 0; 
  adj[2205] = 0; 
  adj[2206] = 0; 
  adj[2207] = 0; 
  adj[2208] = 0; 
  adj[2209] = 1; 
  adj[2210] = 0; 
  adj[2211] = 1; 
  adj[2212] = 0; 
  adj[2213] = 0; 
  adj[2214] = 0; 
  adj[2215] = 0; 
  adj[2216] = 0; 
  adj[2217] = 0; 
  adj[2218] = 0; 
  adj[2219] = 0; 
  adj[2220] = 0; 
  adj[2221] = 0; 
  adj[2222] = 0; 
  adj[2223] = 0; 
  adj[2224] = 0; 
  adj[2225] = 0; 
  adj[2226] = 0; 
  adj[2227] = 0; 
  adj[2228] = 0; 
  adj[2229] = 0; 
  adj[2230] = 0; 
  adj[2231] = 0; 
  adj[2232] = 0; 
  adj[2233] = 0; 
  adj[2234] = 0; 
  adj[2235] = 0; 
  adj[2236] = 0; 
  adj[2237] = 0; 
  adj[2238] = 0; 
  adj[2239] = 0; 
  adj[2240] = 0; 
  adj[2241] = 0; 
  adj[2242] = 0; 
  adj[2243] = 0; 
  adj[2244] = 0; 
  adj[2245] = 0; 
  adj[2246] = 0; 
  adj[2247] = 0; 
  adj[2248] = 0; 
  adj[2249] = 0; 
  adj[2250] = 0; 
  adj[2251] = 0; 
  adj[2252] = 0; 
  adj[2253] = 0; 
  adj[2254] = 0; 
  adj[2255] = 0; 
  adj[2256] = 0; 
  adj[2257] = 0; 
  adj[2258] = 0; 
  adj[2259] = 0; 
  adj[2260] = 0; 
  adj[2261] = 0; 
  adj[2262] = 0; 
  adj[2263] = 0; 
  adj[2264] = 0; 
  adj[2265] = 0; 
  adj[2266] = 0; 
  adj[2267] = 0; 
  adj[2268] = 0; 
  adj[2269] = 0; 
  adj[2270] = 0; 
  adj[2271] = 0; 
  adj[2272] = 0; 
  adj[2273] = 0; 
  adj[2274] = 1; 
  adj[2275] = 0; 
  adj[2276] = 1; 
  adj[2277] = 0; 
  adj[2278] = 0; 
  adj[2279] = 0; 
  adj[2280] = 0; 
  adj[2281] = 0; 
  adj[2282] = 0; 
  adj[2283] = 0; 
  adj[2284] = 0; 
  adj[2285] = 0; 
  adj[2286] = 0; 
  adj[2287] = 0; 
  adj[2288] = 0; 
  adj[2289] = 0; 
  adj[2290] = 0; 
  adj[2291] = 0; 
  adj[2292] = 0; 
  adj[2293] = 0; 
  adj[2294] = 0; 
  adj[2295] = 0; 
  adj[2296] = 0; 
  adj[2297] = 0; 
  adj[2298] = 0; 
  adj[2299] = 0; 
  adj[2300] = 0; 
  adj[2301] = 0; 
  adj[2302] = 0; 
  adj[2303] = 0; 
  adj[2304] = 0; 
  adj[2305] = 0; 
  adj[2306] = 0; 
  adj[2307] = 0; 
  adj[2308] = 0; 
  adj[2309] = 0; 
  adj[2310] = 0; 
  adj[2311] = 0; 
  adj[2312] = 0; 
  adj[2313] = 0; 
  adj[2314] = 0; 
  adj[2315] = 0; 
  adj[2316] = 0; 
  adj[2317] = 0; 
  adj[2318] = 0; 
  adj[2319] = 0; 
  adj[2320] = 0; 
  adj[2321] = 0; 
  adj[2322] = 0; 
  adj[2323] = 0; 
  adj[2324] = 0; 
  adj[2325] = 0; 
  adj[2326] = 0; 
  adj[2327] = 0; 
  adj[2328] = 0; 
  adj[2329] = 0; 
  adj[2330] = 0; 
  adj[2331] = 0; 
  adj[2332] = 0; 
  adj[2333] = 0; 
  adj[2334] = 0; 
  adj[2335] = 0; 
  adj[2336] = 0; 
  adj[2337] = 0; 
  adj[2338] = 0; 
  adj[2339] = 1; 
  adj[2340] = 0; 
  adj[2341] = 1; 
  adj[2342] = 0; 
  adj[2343] = 0; 
  adj[2344] = 0; 
  adj[2345] = 0; 
  adj[2346] = 0; 
  adj[2347] = 0; 
  adj[2348] = 0; 
  adj[2349] = 0; 
  adj[2350] = 0; 
  adj[2351] = 0; 
  adj[2352] = 0; 
  adj[2353] = 0; 
  adj[2354] = 0; 
  adj[2355] = 0; 
  adj[2356] = 0; 
  adj[2357] = 0; 
  adj[2358] = 0; 
  adj[2359] = 0; 
  adj[2360] = 0; 
  adj[2361] = 0; 
  adj[2362] = 0; 
  adj[2363] = 0; 
  adj[2364] = 0; 
  adj[2365] = 0; 
  adj[2366] = 0; 
  adj[2367] = 0; 
  adj[2368] = 0; 
  adj[2369] = 0; 
  adj[2370] = 0; 
  adj[2371] = 0; 
  adj[2372] = 0; 
  adj[2373] = 0; 
  adj[2374] = 0; 
  adj[2375] = 0; 
  adj[2376] = 0; 
  adj[2377] = 0; 
  adj[2378] = 0; 
  adj[2379] = 0; 
  adj[2380] = 0; 
  adj[2381] = 0; 
  adj[2382] = 0; 
  adj[2383] = 0; 
  adj[2384] = 0; 
  adj[2385] = 0; 
  adj[2386] = 0; 
  adj[2387] = 0; 
  adj[2388] = 0; 
  adj[2389] = 0; 
  adj[2390] = 0; 
  adj[2391] = 0; 
  adj[2392] = 0; 
  adj[2393] = 0; 
  adj[2394] = 0; 
  adj[2395] = 0; 
  adj[2396] = 0; 
  adj[2397] = 0; 
  adj[2398] = 0; 
  adj[2399] = 0; 
  adj[2400] = 0; 
  adj[2401] = 0; 
  adj[2402] = 0; 
  adj[2403] = 0; 
  adj[2404] = 1; 
  adj[2405] = 0; 
  adj[2406] = 1; 
  adj[2407] = 0; 
  adj[2408] = 0; 
  adj[2409] = 0; 
  adj[2410] = 0; 
  adj[2411] = 0; 
  adj[2412] = 0; 
  adj[2413] = 0; 
  adj[2414] = 0; 
  adj[2415] = 0; 
  adj[2416] = 0; 
  adj[2417] = 0; 
  adj[2418] = 0; 
  adj[2419] = 0; 
  adj[2420] = 0; 
  adj[2421] = 0; 
  adj[2422] = 0; 
  adj[2423] = 0; 
  adj[2424] = 0; 
  adj[2425] = 0; 
  adj[2426] = 0; 
  adj[2427] = 0; 
  adj[2428] = 0; 
  adj[2429] = 0; 
  adj[2430] = 0; 
  adj[2431] = 0; 
  adj[2432] = 0; 
  adj[2433] = 0; 
  adj[2434] = 0; 
  adj[2435] = 0; 
  adj[2436] = 0; 
  adj[2437] = 0; 
  adj[2438] = 0; 
  adj[2439] = 0; 
  adj[2440] = 0; 
  adj[2441] = 0; 
  adj[2442] = 0; 
  adj[2443] = 0; 
  adj[2444] = 0; 
  adj[2445] = 0; 
  adj[2446] = 0; 
  adj[2447] = 0; 
  adj[2448] = 0; 
  adj[2449] = 0; 
  adj[2450] = 0; 
  adj[2451] = 0; 
  adj[2452] = 0; 
  adj[2453] = 0; 
  adj[2454] = 0; 
  adj[2455] = 0; 
  adj[2456] = 0; 
  adj[2457] = 0; 
  adj[2458] = 0; 
  adj[2459] = 0; 
  adj[2460] = 0; 
  adj[2461] = 0; 
  adj[2462] = 0; 
  adj[2463] = 0; 
  adj[2464] = 0; 
  adj[2465] = 0; 
  adj[2466] = 0; 
  adj[2467] = 0; 
  adj[2468] = 0; 
  adj[2469] = 1; 
  adj[2470] = 0; 
  adj[2471] = 1; 
  adj[2472] = 0; 
  adj[2473] = 0; 
  adj[2474] = 0; 
  adj[2475] = 0; 
  adj[2476] = 0; 
  adj[2477] = 0; 
  adj[2478] = 0; 
  adj[2479] = 0; 
  adj[2480] = 0; 
  adj[2481] = 0; 
  adj[2482] = 0; 
  adj[2483] = 0; 
  adj[2484] = 0; 
  adj[2485] = 0; 
  adj[2486] = 0; 
  adj[2487] = 0; 
  adj[2488] = 0; 
  adj[2489] = 0; 
  adj[2490] = 0; 
  adj[2491] = 0; 
  adj[2492] = 0; 
  adj[2493] = 0; 
  adj[2494] = 0; 
  adj[2495] = 0; 
  adj[2496] = 0; 
  adj[2497] = 0; 
  adj[2498] = 0; 
  adj[2499] = 0; 
  adj[2500] = 0; 
  adj[2501] = 0; 
  adj[2502] = 0; 
  adj[2503] = 0; 
  adj[2504] = 0; 
  adj[2505] = 0; 
  adj[2506] = 0; 
  adj[2507] = 0; 
  adj[2508] = 0; 
  adj[2509] = 0; 
  adj[2510] = 0; 
  adj[2511] = 0; 
  adj[2512] = 0; 
  adj[2513] = 0; 
  adj[2514] = 0; 
  adj[2515] = 0; 
  adj[2516] = 0; 
  adj[2517] = 0; 
  adj[2518] = 0; 
  adj[2519] = 0; 
  adj[2520] = 0; 
  adj[2521] = 0; 
  adj[2522] = 0; 
  adj[2523] = 1; 
  adj[2524] = 0; 
  adj[2525] = 0; 
  adj[2526] = 0; 
  adj[2527] = 0; 
  adj[2528] = 0; 
  adj[2529] = 0; 
  adj[2530] = 0; 
  adj[2531] = 0; 
  adj[2532] = 0; 
  adj[2533] = 0; 
  adj[2534] = 1; 
  adj[2535] = 0; 
  adj[2536] = 1; 
  adj[2537] = 0; 
  adj[2538] = 0; 
  adj[2539] = 0; 
  adj[2540] = 0; 
  adj[2541] = 0; 
  adj[2542] = 0; 
  adj[2543] = 0; 
  adj[2544] = 0; 
  adj[2545] = 0; 
  adj[2546] = 0; 
  adj[2547] = 0; 
  adj[2548] = 0; 
  adj[2549] = 0; 
  adj[2550] = 0; 
  adj[2551] = 0; 
  adj[2552] = 0; 
  adj[2553] = 0; 
  adj[2554] = 0; 
  adj[2555] = 0; 
  adj[2556] = 0; 
  adj[2557] = 0; 
  adj[2558] = 0; 
  adj[2559] = 0; 
  adj[2560] = 0; 
  adj[2561] = 0; 
  adj[2562] = 0; 
  adj[2563] = 0; 
  adj[2564] = 0; 
  adj[2565] = 0; 
  adj[2566] = 0; 
  adj[2567] = 0; 
  adj[2568] = 0; 
  adj[2569] = 0; 
  adj[2570] = 0; 
  adj[2571] = 0; 
  adj[2572] = 0; 
  adj[2573] = 0; 
  adj[2574] = 0; 
  adj[2575] = 0; 
  adj[2576] = 0; 
  adj[2577] = 0; 
  adj[2578] = 0; 
  adj[2579] = 0; 
  adj[2580] = 0; 
  adj[2581] = 0; 
  adj[2582] = 0; 
  adj[2583] = 0; 
  adj[2584] = 0; 
  adj[2585] = 0; 
  adj[2586] = 0; 
  adj[2587] = 0; 
  adj[2588] = 0; 
  adj[2589] = 0; 
  adj[2590] = 0; 
  adj[2591] = 0; 
  adj[2592] = 0; 
  adj[2593] = 0; 
  adj[2594] = 0; 
  adj[2595] = 0; 
  adj[2596] = 0; 
  adj[2597] = 0; 
  adj[2598] = 0; 
  adj[2599] = 1; 
  adj[2600] = 0; 
  adj[2601] = 1; 
  adj[2602] = 0; 
  adj[2603] = 0; 
  adj[2604] = 0; 
  adj[2605] = 0; 
  adj[2606] = 0; 
  adj[2607] = 0; 
  adj[2608] = 0; 
  adj[2609] = 0; 
  adj[2610] = 0; 
  adj[2611] = 0; 
  adj[2612] = 0; 
  adj[2613] = 0; 
  adj[2614] = 0; 
  adj[2615] = 0; 
  adj[2616] = 0; 
  adj[2617] = 0; 
  adj[2618] = 0; 
  adj[2619] = 0; 
  adj[2620] = 0; 
  adj[2621] = 0; 
  adj[2622] = 0; 
  adj[2623] = 0; 
  adj[2624] = 0; 
  adj[2625] = 0; 
  adj[2626] = 0; 
  adj[2627] = 0; 
  adj[2628] = 0; 
  adj[2629] = 0; 
  adj[2630] = 0; 
  adj[2631] = 0; 
  adj[2632] = 0; 
  adj[2633] = 0; 
  adj[2634] = 0; 
  adj[2635] = 0; 
  adj[2636] = 0; 
  adj[2637] = 0; 
  adj[2638] = 0; 
  adj[2639] = 0; 
  adj[2640] = 0; 
  adj[2641] = 0; 
  adj[2642] = 0; 
  adj[2643] = 0; 
  adj[2644] = 0; 
  adj[2645] = 0; 
  adj[2646] = 0; 
  adj[2647] = 0; 
  adj[2648] = 0; 
  adj[2649] = 0; 
  adj[2650] = 0; 
  adj[2651] = 0; 
  adj[2652] = 0; 
  adj[2653] = 0; 
  adj[2654] = 0; 
  adj[2655] = 0; 
  adj[2656] = 0; 
  adj[2657] = 0; 
  adj[2658] = 0; 
  adj[2659] = 0; 
  adj[2660] = 0; 
  adj[2661] = 0; 
  adj[2662] = 0; 
  adj[2663] = 0; 
  adj[2664] = 1; 
  adj[2665] = 0; 
  adj[2666] = 1; 
  adj[2667] = 0; 
  adj[2668] = 0; 
  adj[2669] = 0; 
  adj[2670] = 0; 
  adj[2671] = 0; 
  adj[2672] = 0; 
  adj[2673] = 0; 
  adj[2674] = 0; 
  adj[2675] = 0; 
  adj[2676] = 0; 
  adj[2677] = 0; 
  adj[2678] = 0; 
  adj[2679] = 0; 
  adj[2680] = 0; 
  adj[2681] = 0; 
  adj[2682] = 0; 
  adj[2683] = 0; 
  adj[2684] = 0; 
  adj[2685] = 0; 
  adj[2686] = 0; 
  adj[2687] = 0; 
  adj[2688] = 0; 
  adj[2689] = 0; 
  adj[2690] = 0; 
  adj[2691] = 0; 
  adj[2692] = 0; 
  adj[2693] = 0; 
  adj[2694] = 0; 
  adj[2695] = 0; 
  adj[2696] = 0; 
  adj[2697] = 0; 
  adj[2698] = 0; 
  adj[2699] = 0; 
  adj[2700] = 0; 
  adj[2701] = 0; 
  adj[2702] = 0; 
  adj[2703] = 0; 
  adj[2704] = 0; 
  adj[2705] = 0; 
  adj[2706] = 0; 
  adj[2707] = 0; 
  adj[2708] = 0; 
  adj[2709] = 0; 
  adj[2710] = 0; 
  adj[2711] = 0; 
  adj[2712] = 0; 
  adj[2713] = 0; 
  adj[2714] = 0; 
  adj[2715] = 0; 
  adj[2716] = 0; 
  adj[2717] = 0; 
  adj[2718] = 0; 
  adj[2719] = 0; 
  adj[2720] = 0; 
  adj[2721] = 0; 
  adj[2722] = 0; 
  adj[2723] = 0; 
  adj[2724] = 0; 
  adj[2725] = 0; 
  adj[2726] = 0; 
  adj[2727] = 0; 
  adj[2728] = 0; 
  adj[2729] = 1; 
  adj[2730] = 0; 
  adj[2731] = 1; 
  adj[2732] = 0; 
  adj[2733] = 0; 
  adj[2734] = 0; 
  adj[2735] = 0; 
  adj[2736] = 0; 
  adj[2737] = 0; 
  adj[2738] = 0; 
  adj[2739] = 0; 
  adj[2740] = 0; 
  adj[2741] = 0; 
  adj[2742] = 0; 
  adj[2743] = 0; 
  adj[2744] = 0; 
  adj[2745] = 0; 
  adj[2746] = 0; 
  adj[2747] = 0; 
  adj[2748] = 0; 
  adj[2749] = 0; 
  adj[2750] = 0; 
  adj[2751] = 0; 
  adj[2752] = 0; 
  adj[2753] = 0; 
  adj[2754] = 0; 
  adj[2755] = 0; 
  adj[2756] = 0; 
  adj[2757] = 0; 
  adj[2758] = 0; 
  adj[2759] = 0; 
  adj[2760] = 0; 
  adj[2761] = 0; 
  adj[2762] = 0; 
  adj[2763] = 0; 
  adj[2764] = 0; 
  adj[2765] = 0; 
  adj[2766] = 0; 
  adj[2767] = 0; 
  adj[2768] = 0; 
  adj[2769] = 0; 
  adj[2770] = 0; 
  adj[2771] = 0; 
  adj[2772] = 0; 
  adj[2773] = 0; 
  adj[2774] = 0; 
  adj[2775] = 0; 
  adj[2776] = 0; 
  adj[2777] = 0; 
  adj[2778] = 0; 
  adj[2779] = 0; 
  adj[2780] = 0; 
  adj[2781] = 0; 
  adj[2782] = 0; 
  adj[2783] = 0; 
  adj[2784] = 0; 
  adj[2785] = 0; 
  adj[2786] = 0; 
  adj[2787] = 0; 
  adj[2788] = 0; 
  adj[2789] = 0; 
  adj[2790] = 0; 
  adj[2791] = 0; 
  adj[2792] = 0; 
  adj[2793] = 0; 
  adj[2794] = 1; 
  adj[2795] = 0; 
  adj[2796] = 1; 
  adj[2797] = 0; 
  adj[2798] = 0; 
  adj[2799] = 0; 
  adj[2800] = 0; 
  adj[2801] = 0; 
  adj[2802] = 0; 
  adj[2803] = 0; 
  adj[2804] = 0; 
  adj[2805] = 0; 
  adj[2806] = 0; 
  adj[2807] = 0; 
  adj[2808] = 0; 
  adj[2809] = 0; 
  adj[2810] = 0; 
  adj[2811] = 0; 
  adj[2812] = 0; 
  adj[2813] = 0; 
  adj[2814] = 0; 
  adj[2815] = 0; 
  adj[2816] = 0; 
  adj[2817] = 0; 
  adj[2818] = 0; 
  adj[2819] = 0; 
  adj[2820] = 0; 
  adj[2821] = 0; 
  adj[2822] = 0; 
  adj[2823] = 0; 
  adj[2824] = 0; 
  adj[2825] = 0; 
  adj[2826] = 0; 
  adj[2827] = 0; 
  adj[2828] = 0; 
  adj[2829] = 0; 
  adj[2830] = 0; 
  adj[2831] = 0; 
  adj[2832] = 0; 
  adj[2833] = 0; 
  adj[2834] = 0; 
  adj[2835] = 0; 
  adj[2836] = 0; 
  adj[2837] = 0; 
  adj[2838] = 0; 
  adj[2839] = 0; 
  adj[2840] = 0; 
  adj[2841] = 0; 
  adj[2842] = 0; 
  adj[2843] = 0; 
  adj[2844] = 0; 
  adj[2845] = 0; 
  adj[2846] = 0; 
  adj[2847] = 0; 
  adj[2848] = 0; 
  adj[2849] = 0; 
  adj[2850] = 0; 
  adj[2851] = 0; 
  adj[2852] = 0; 
  adj[2853] = 0; 
  adj[2854] = 0; 
  adj[2855] = 0; 
  adj[2856] = 0; 
  adj[2857] = 0; 
  adj[2858] = 0; 
  adj[2859] = 1; 
  adj[2860] = 0; 
  adj[2861] = 1; 
  adj[2862] = 0; 
  adj[2863] = 0; 
  adj[2864] = 0; 
  adj[2865] = 0; 
  adj[2866] = 0; 
  adj[2867] = 0; 
  adj[2868] = 0; 
  adj[2869] = 0; 
  adj[2870] = 0; 
  adj[2871] = 0; 
  adj[2872] = 0; 
  adj[2873] = 0; 
  adj[2874] = 0; 
  adj[2875] = 0; 
  adj[2876] = 0; 
  adj[2877] = 0; 
  adj[2878] = 0; 
  adj[2879] = 0; 
  adj[2880] = 0; 
  adj[2881] = 0; 
  adj[2882] = 0; 
  adj[2883] = 0; 
  adj[2884] = 0; 
  adj[2885] = 0; 
  adj[2886] = 0; 
  adj[2887] = 0; 
  adj[2888] = 0; 
  adj[2889] = 0; 
  adj[2890] = 0; 
  adj[2891] = 0; 
  adj[2892] = 0; 
  adj[2893] = 0; 
  adj[2894] = 0; 
  adj[2895] = 0; 
  adj[2896] = 0; 
  adj[2897] = 0; 
  adj[2898] = 0; 
  adj[2899] = 0; 
  adj[2900] = 0; 
  adj[2901] = 0; 
  adj[2902] = 0; 
  adj[2903] = 0; 
  adj[2904] = 0; 
  adj[2905] = 0; 
  adj[2906] = 0; 
  adj[2907] = 0; 
  adj[2908] = 0; 
  adj[2909] = 0; 
  adj[2910] = 0; 
  adj[2911] = 0; 
  adj[2912] = 0; 
  adj[2913] = 0; 
  adj[2914] = 0; 
  adj[2915] = 0; 
  adj[2916] = 0; 
  adj[2917] = 0; 
  adj[2918] = 0; 
  adj[2919] = 0; 
  adj[2920] = 0; 
  adj[2921] = 0; 
  adj[2922] = 0; 
  adj[2923] = 0; 
  adj[2924] = 1; 
  adj[2925] = 0; 
  adj[2926] = 1; 
  adj[2927] = 0; 
  adj[2928] = 0; 
  adj[2929] = 0; 
  adj[2930] = 0; 
  adj[2931] = 0; 
  adj[2932] = 0; 
  adj[2933] = 0; 
  adj[2934] = 0; 
  adj[2935] = 0; 
  adj[2936] = 0; 
  adj[2937] = 0; 
  adj[2938] = 0; 
  adj[2939] = 0; 
  adj[2940] = 0; 
  adj[2941] = 0; 
  adj[2942] = 0; 
  adj[2943] = 0; 
  adj[2944] = 0; 
  adj[2945] = 0; 
  adj[2946] = 0; 
  adj[2947] = 0; 
  adj[2948] = 0; 
  adj[2949] = 0; 
  adj[2950] = 0; 
  adj[2951] = 0; 
  adj[2952] = 0; 
  adj[2953] = 0; 
  adj[2954] = 0; 
  adj[2955] = 0; 
  adj[2956] = 0; 
  adj[2957] = 0; 
  adj[2958] = 0; 
  adj[2959] = 0; 
  adj[2960] = 0; 
  adj[2961] = 0; 
  adj[2962] = 0; 
  adj[2963] = 0; 
  adj[2964] = 0; 
  adj[2965] = 0; 
  adj[2966] = 0; 
  adj[2967] = 0; 
  adj[2968] = 0; 
  adj[2969] = 0; 
  adj[2970] = 0; 
  adj[2971] = 0; 
  adj[2972] = 0; 
  adj[2973] = 0; 
  adj[2974] = 0; 
  adj[2975] = 0; 
  adj[2976] = 0; 
  adj[2977] = 0; 
  adj[2978] = 0; 
  adj[2979] = 0; 
  adj[2980] = 0; 
  adj[2981] = 0; 
  adj[2982] = 0; 
  adj[2983] = 0; 
  adj[2984] = 0; 
  adj[2985] = 0; 
  adj[2986] = 0; 
  adj[2987] = 0; 
  adj[2988] = 0; 
  adj[2989] = 1; 
  adj[2990] = 0; 
  adj[2991] = 1; 
  adj[2992] = 0; 
  adj[2993] = 0; 
  adj[2994] = 0; 
  adj[2995] = 0; 
  adj[2996] = 0; 
  adj[2997] = 0; 
  adj[2998] = 0; 
  adj[2999] = 0; 
  adj[3000] = 0; 
  adj[3001] = 0; 
  adj[3002] = 0; 
  adj[3003] = 0; 
  adj[3004] = 0; 
  adj[3005] = 0; 
  adj[3006] = 0; 
  adj[3007] = 0; 
  adj[3008] = 0; 
  adj[3009] = 0; 
  adj[3010] = 0; 
  adj[3011] = 0; 
  adj[3012] = 0; 
  adj[3013] = 0; 
  adj[3014] = 0; 
  adj[3015] = 0; 
  adj[3016] = 0; 
  adj[3017] = 0; 
  adj[3018] = 0; 
  adj[3019] = 0; 
  adj[3020] = 0; 
  adj[3021] = 0; 
  adj[3022] = 0; 
  adj[3023] = 0; 
  adj[3024] = 0; 
  adj[3025] = 0; 
  adj[3026] = 0; 
  adj[3027] = 0; 
  adj[3028] = 0; 
  adj[3029] = 0; 
  adj[3030] = 0; 
  adj[3031] = 0; 
  adj[3032] = 0; 
  adj[3033] = 0; 
  adj[3034] = 0; 
  adj[3035] = 0; 
  adj[3036] = 0; 
  adj[3037] = 0; 
  adj[3038] = 0; 
  adj[3039] = 0; 
  adj[3040] = 0; 
  adj[3041] = 0; 
  adj[3042] = 0; 
  adj[3043] = 0; 
  adj[3044] = 0; 
  adj[3045] = 0; 
  adj[3046] = 0; 
  adj[3047] = 0; 
  adj[3048] = 0; 
  adj[3049] = 0; 
  adj[3050] = 0; 
  adj[3051] = 0; 
  adj[3052] = 0; 
  adj[3053] = 0; 
  adj[3054] = 1; 
  adj[3055] = 0; 
  adj[3056] = 1; 
  adj[3057] = 0; 
  adj[3058] = 0; 
  adj[3059] = 0; 
  adj[3060] = 0; 
  adj[3061] = 0; 
  adj[3062] = 0; 
  adj[3063] = 0; 
  adj[3064] = 0; 
  adj[3065] = 0; 
  adj[3066] = 0; 
  adj[3067] = 0; 
  adj[3068] = 0; 
  adj[3069] = 0; 
  adj[3070] = 0; 
  adj[3071] = 0; 
  adj[3072] = 0; 
  adj[3073] = 0; 
  adj[3074] = 0; 
  adj[3075] = 0; 
  adj[3076] = 0; 
  adj[3077] = 0; 
  adj[3078] = 0; 
  adj[3079] = 0; 
  adj[3080] = 0; 
  adj[3081] = 0; 
  adj[3082] = 0; 
  adj[3083] = 0; 
  adj[3084] = 0; 
  adj[3085] = 0; 
  adj[3086] = 0; 
  adj[3087] = 0; 
  adj[3088] = 0; 
  adj[3089] = 0; 
  adj[3090] = 0; 
  adj[3091] = 0; 
  adj[3092] = 0; 
  adj[3093] = 0; 
  adj[3094] = 0; 
  adj[3095] = 0; 
  adj[3096] = 0; 
  adj[3097] = 0; 
  adj[3098] = 0; 
  adj[3099] = 0; 
  adj[3100] = 0; 
  adj[3101] = 0; 
  adj[3102] = 0; 
  adj[3103] = 0; 
  adj[3104] = 0; 
  adj[3105] = 0; 
  adj[3106] = 0; 
  adj[3107] = 0; 
  adj[3108] = 0; 
  adj[3109] = 0; 
  adj[3110] = 0; 
  adj[3111] = 0; 
  adj[3112] = 0; 
  adj[3113] = 0; 
  adj[3114] = 0; 
  adj[3115] = 0; 
  adj[3116] = 0; 
  adj[3117] = 0; 
  adj[3118] = 0; 
  adj[3119] = 1; 
  adj[3120] = 0; 
  adj[3121] = 1; 
  adj[3122] = 0; 
  adj[3123] = 0; 
  adj[3124] = 0; 
  adj[3125] = 0; 
  adj[3126] = 0; 
  adj[3127] = 0; 
  adj[3128] = 0; 
  adj[3129] = 0; 
  adj[3130] = 0; 
  adj[3131] = 0; 
  adj[3132] = 0; 
  adj[3133] = 0; 
  adj[3134] = 0; 
  adj[3135] = 0; 
  adj[3136] = 0; 
  adj[3137] = 0; 
  adj[3138] = 0; 
  adj[3139] = 0; 
  adj[3140] = 0; 
  adj[3141] = 0; 
  adj[3142] = 0; 
  adj[3143] = 0; 
  adj[3144] = 0; 
  adj[3145] = 0; 
  adj[3146] = 0; 
  adj[3147] = 0; 
  adj[3148] = 0; 
  adj[3149] = 0; 
  adj[3150] = 0; 
  adj[3151] = 0; 
  adj[3152] = 0; 
  adj[3153] = 0; 
  adj[3154] = 0; 
  adj[3155] = 0; 
  adj[3156] = 0; 
  adj[3157] = 0; 
  adj[3158] = 0; 
  adj[3159] = 0; 
  adj[3160] = 0; 
  adj[3161] = 0; 
  adj[3162] = 0; 
  adj[3163] = 0; 
  adj[3164] = 0; 
  adj[3165] = 0; 
  adj[3166] = 0; 
  adj[3167] = 0; 
  adj[3168] = 0; 
  adj[3169] = 0; 
  adj[3170] = 0; 
  adj[3171] = 0; 
  adj[3172] = 0; 
  adj[3173] = 0; 
  adj[3174] = 0; 
  adj[3175] = 0; 
  adj[3176] = 0; 
  adj[3177] = 0; 
  adj[3178] = 0; 
  adj[3179] = 0; 
  adj[3180] = 0; 
  adj[3181] = 0; 
  adj[3182] = 0; 
  adj[3183] = 0; 
  adj[3184] = 1; 
  adj[3185] = 0; 
  adj[3186] = 1; 
  adj[3187] = 0; 
  adj[3188] = 0; 
  adj[3189] = 0; 
  adj[3190] = 0; 
  adj[3191] = 0; 
  adj[3192] = 0; 
  adj[3193] = 0; 
  adj[3194] = 0; 
  adj[3195] = 0; 
  adj[3196] = 0; 
  adj[3197] = 0; 
  adj[3198] = 0; 
  adj[3199] = 0; 
  adj[3200] = 0; 
  adj[3201] = 0; 
  adj[3202] = 0; 
  adj[3203] = 0; 
  adj[3204] = 0; 
  adj[3205] = 0; 
  adj[3206] = 0; 
  adj[3207] = 0; 
  adj[3208] = 0; 
  adj[3209] = 0; 
  adj[3210] = 0; 
  adj[3211] = 0; 
  adj[3212] = 0; 
  adj[3213] = 0; 
  adj[3214] = 0; 
  adj[3215] = 0; 
  adj[3216] = 0; 
  adj[3217] = 0; 
  adj[3218] = 0; 
  adj[3219] = 0; 
  adj[3220] = 0; 
  adj[3221] = 0; 
  adj[3222] = 0; 
  adj[3223] = 0; 
  adj[3224] = 0; 
  adj[3225] = 0; 
  adj[3226] = 0; 
  adj[3227] = 0; 
  adj[3228] = 0; 
  adj[3229] = 0; 
  adj[3230] = 0; 
  adj[3231] = 0; 
  adj[3232] = 0; 
  adj[3233] = 0; 
  adj[3234] = 0; 
  adj[3235] = 0; 
  adj[3236] = 0; 
  adj[3237] = 0; 
  adj[3238] = 0; 
  adj[3239] = 0; 
  adj[3240] = 0; 
  adj[3241] = 0; 
  adj[3242] = 0; 
  adj[3243] = 0; 
  adj[3244] = 0; 
  adj[3245] = 0; 
  adj[3246] = 0; 
  adj[3247] = 0; 
  adj[3248] = 0; 
  adj[3249] = 1; 
  adj[3250] = 0; 
  adj[3251] = 1; 
  adj[3252] = 0; 
  adj[3253] = 0; 
  adj[3254] = 0; 
  adj[3255] = 0; 
  adj[3256] = 0; 
  adj[3257] = 0; 
  adj[3258] = 0; 
  adj[3259] = 0; 
  adj[3260] = 0; 
  adj[3261] = 0; 
  adj[3262] = 0; 
  adj[3263] = 0; 
  adj[3264] = 0; 
  adj[3265] = 0; 
  adj[3266] = 0; 
  adj[3267] = 0; 
  adj[3268] = 0; 
  adj[3269] = 0; 
  adj[3270] = 0; 
  adj[3271] = 0; 
  adj[3272] = 0; 
  adj[3273] = 0; 
  adj[3274] = 0; 
  adj[3275] = 0; 
  adj[3276] = 0; 
  adj[3277] = 0; 
  adj[3278] = 0; 
  adj[3279] = 0; 
  adj[3280] = 0; 
  adj[3281] = 0; 
  adj[3282] = 0; 
  adj[3283] = 0; 
  adj[3284] = 0; 
  adj[3285] = 0; 
  adj[3286] = 0; 
  adj[3287] = 0; 
  adj[3288] = 0; 
  adj[3289] = 0; 
  adj[3290] = 0; 
  adj[3291] = 0; 
  adj[3292] = 0; 
  adj[3293] = 0; 
  adj[3294] = 0; 
  adj[3295] = 0; 
  adj[3296] = 0; 
  adj[3297] = 0; 
  adj[3298] = 0; 
  adj[3299] = 0; 
  adj[3300] = 0; 
  adj[3301] = 0; 
  adj[3302] = 0; 
  adj[3303] = 0; 
  adj[3304] = 0; 
  adj[3305] = 0; 
  adj[3306] = 0; 
  adj[3307] = 0; 
  adj[3308] = 0; 
  adj[3309] = 0; 
  adj[3310] = 0; 
  adj[3311] = 0; 
  adj[3312] = 0; 
  adj[3313] = 0; 
  adj[3314] = 1; 
  adj[3315] = 0; 
  adj[3316] = 1; 
  adj[3317] = 0; 
  adj[3318] = 0; 
  adj[3319] = 0; 
  adj[3320] = 0; 
  adj[3321] = 0; 
  adj[3322] = 0; 
  adj[3323] = 0; 
  adj[3324] = 0; 
  adj[3325] = 0; 
  adj[3326] = 0; 
  adj[3327] = 0; 
  adj[3328] = 0; 
  adj[3329] = 0; 
  adj[3330] = 0; 
  adj[3331] = 0; 
  adj[3332] = 0; 
  adj[3333] = 0; 
  adj[3334] = 0; 
  adj[3335] = 0; 
  adj[3336] = 0; 
  adj[3337] = 0; 
  adj[3338] = 0; 
  adj[3339] = 0; 
  adj[3340] = 0; 
  adj[3341] = 0; 
  adj[3342] = 0; 
  adj[3343] = 0; 
  adj[3344] = 0; 
  adj[3345] = 1; 
  adj[3346] = 0; 
  adj[3347] = 0; 
  adj[3348] = 0; 
  adj[3349] = 0; 
  adj[3350] = 0; 
  adj[3351] = 0; 
  adj[3352] = 0; 
  adj[3353] = 0; 
  adj[3354] = 0; 
  adj[3355] = 0; 
  adj[3356] = 0; 
  adj[3357] = 0; 
  adj[3358] = 0; 
  adj[3359] = 0; 
  adj[3360] = 0; 
  adj[3361] = 0; 
  adj[3362] = 0; 
  adj[3363] = 0; 
  adj[3364] = 0; 
  adj[3365] = 0; 
  adj[3366] = 0; 
  adj[3367] = 0; 
  adj[3368] = 0; 
  adj[3369] = 0; 
  adj[3370] = 0; 
  adj[3371] = 0; 
  adj[3372] = 0; 
  adj[3373] = 0; 
  adj[3374] = 0; 
  adj[3375] = 0; 
  adj[3376] = 0; 
  adj[3377] = 0; 
  adj[3378] = 0; 
  adj[3379] = 1; 
  adj[3380] = 0; 
  adj[3381] = 1; 
  adj[3382] = 0; 
  adj[3383] = 0; 
  adj[3384] = 0; 
  adj[3385] = 0; 
  adj[3386] = 0; 
  adj[3387] = 0; 
  adj[3388] = 0; 
  adj[3389] = 0; 
  adj[3390] = 0; 
  adj[3391] = 0; 
  adj[3392] = 0; 
  adj[3393] = 0; 
  adj[3394] = 0; 
  adj[3395] = 0; 
  adj[3396] = 0; 
  adj[3397] = 0; 
  adj[3398] = 0; 
  adj[3399] = 0; 
  adj[3400] = 0; 
  adj[3401] = 0; 
  adj[3402] = 0; 
  adj[3403] = 0; 
  adj[3404] = 0; 
  adj[3405] = 0; 
  adj[3406] = 0; 
  adj[3407] = 0; 
  adj[3408] = 0; 
  adj[3409] = 0; 
  adj[3410] = 0; 
  adj[3411] = 0; 
  adj[3412] = 0; 
  adj[3413] = 0; 
  adj[3414] = 0; 
  adj[3415] = 0; 
  adj[3416] = 0; 
  adj[3417] = 0; 
  adj[3418] = 0; 
  adj[3419] = 0; 
  adj[3420] = 0; 
  adj[3421] = 0; 
  adj[3422] = 0; 
  adj[3423] = 0; 
  adj[3424] = 0; 
  adj[3425] = 0; 
  adj[3426] = 0; 
  adj[3427] = 0; 
  adj[3428] = 0; 
  adj[3429] = 0; 
  adj[3430] = 0; 
  adj[3431] = 0; 
  adj[3432] = 0; 
  adj[3433] = 0; 
  adj[3434] = 0; 
  adj[3435] = 0; 
  adj[3436] = 0; 
  adj[3437] = 0; 
  adj[3438] = 0; 
  adj[3439] = 0; 
  adj[3440] = 0; 
  adj[3441] = 0; 
  adj[3442] = 0; 
  adj[3443] = 0; 
  adj[3444] = 1; 
  adj[3445] = 0; 
  adj[3446] = 1; 
  adj[3447] = 0; 
  adj[3448] = 0; 
  adj[3449] = 0; 
  adj[3450] = 0; 
  adj[3451] = 0; 
  adj[3452] = 0; 
  adj[3453] = 0; 
  adj[3454] = 0; 
  adj[3455] = 0; 
  adj[3456] = 0; 
  adj[3457] = 0; 
  adj[3458] = 0; 
  adj[3459] = 0; 
  adj[3460] = 0; 
  adj[3461] = 0; 
  adj[3462] = 0; 
  adj[3463] = 0; 
  adj[3464] = 0; 
  adj[3465] = 0; 
  adj[3466] = 0; 
  adj[3467] = 0; 
  adj[3468] = 0; 
  adj[3469] = 0; 
  adj[3470] = 0; 
  adj[3471] = 0; 
  adj[3472] = 0; 
  adj[3473] = 0; 
  adj[3474] = 0; 
  adj[3475] = 0; 
  adj[3476] = 0; 
  adj[3477] = 0; 
  adj[3478] = 0; 
  adj[3479] = 0; 
  adj[3480] = 0; 
  adj[3481] = 0; 
  adj[3482] = 0; 
  adj[3483] = 0; 
  adj[3484] = 0; 
  adj[3485] = 0; 
  adj[3486] = 0; 
  adj[3487] = 0; 
  adj[3488] = 0; 
  adj[3489] = 0; 
  adj[3490] = 0; 
  adj[3491] = 0; 
  adj[3492] = 0; 
  adj[3493] = 0; 
  adj[3494] = 0; 
  adj[3495] = 0; 
  adj[3496] = 0; 
  adj[3497] = 0; 
  adj[3498] = 0; 
  adj[3499] = 0; 
  adj[3500] = 0; 
  adj[3501] = 0; 
  adj[3502] = 0; 
  adj[3503] = 0; 
  adj[3504] = 0; 
  adj[3505] = 0; 
  adj[3506] = 0; 
  adj[3507] = 0; 
  adj[3508] = 0; 
  adj[3509] = 1; 
  adj[3510] = 0; 
  adj[3511] = 1; 
  adj[3512] = 0; 
  adj[3513] = 0; 
  adj[3514] = 0; 
  adj[3515] = 0; 
  adj[3516] = 0; 
  adj[3517] = 0; 
  adj[3518] = 0; 
  adj[3519] = 0; 
  adj[3520] = 0; 
  adj[3521] = 0; 
  adj[3522] = 0; 
  adj[3523] = 0; 
  adj[3524] = 0; 
  adj[3525] = 0; 
  adj[3526] = 0; 
  adj[3527] = 0; 
  adj[3528] = 0; 
  adj[3529] = 0; 
  adj[3530] = 0; 
  adj[3531] = 0; 
  adj[3532] = 0; 
  adj[3533] = 0; 
  adj[3534] = 0; 
  adj[3535] = 0; 
  adj[3536] = 0; 
  adj[3537] = 0; 
  adj[3538] = 0; 
  adj[3539] = 0; 
  adj[3540] = 0; 
  adj[3541] = 0; 
  adj[3542] = 0; 
  adj[3543] = 0; 
  adj[3544] = 0; 
  adj[3545] = 0; 
  adj[3546] = 0; 
  adj[3547] = 0; 
  adj[3548] = 0; 
  adj[3549] = 0; 
  adj[3550] = 0; 
  adj[3551] = 0; 
  adj[3552] = 0; 
  adj[3553] = 0; 
  adj[3554] = 0; 
  adj[3555] = 0; 
  adj[3556] = 0; 
  adj[3557] = 0; 
  adj[3558] = 0; 
  adj[3559] = 0; 
  adj[3560] = 0; 
  adj[3561] = 0; 
  adj[3562] = 0; 
  adj[3563] = 0; 
  adj[3564] = 0; 
  adj[3565] = 0; 
  adj[3566] = 0; 
  adj[3567] = 0; 
  adj[3568] = 0; 
  adj[3569] = 0; 
  adj[3570] = 0; 
  adj[3571] = 0; 
  adj[3572] = 0; 
  adj[3573] = 0; 
  adj[3574] = 1; 
  adj[3575] = 0; 
  adj[3576] = 1; 
  adj[3577] = 0; 
  adj[3578] = 0; 
  adj[3579] = 0; 
  adj[3580] = 0; 
  adj[3581] = 0; 
  adj[3582] = 0; 
  adj[3583] = 0; 
  adj[3584] = 0; 
  adj[3585] = 0; 
  adj[3586] = 0; 
  adj[3587] = 0; 
  adj[3588] = 0; 
  adj[3589] = 0; 
  adj[3590] = 0; 
  adj[3591] = 0; 
  adj[3592] = 0; 
  adj[3593] = 0; 
  adj[3594] = 0; 
  adj[3595] = 0; 
  adj[3596] = 0; 
  adj[3597] = 0; 
  adj[3598] = 0; 
  adj[3599] = 0; 
  adj[3600] = 0; 
  adj[3601] = 0; 
  adj[3602] = 0; 
  adj[3603] = 0; 
  adj[3604] = 0; 
  adj[3605] = 0; 
  adj[3606] = 0; 
  adj[3607] = 0; 
  adj[3608] = 0; 
  adj[3609] = 0; 
  adj[3610] = 0; 
  adj[3611] = 0; 
  adj[3612] = 0; 
  adj[3613] = 0; 
  adj[3614] = 0; 
  adj[3615] = 0; 
  adj[3616] = 0; 
  adj[3617] = 0; 
  adj[3618] = 0; 
  adj[3619] = 0; 
  adj[3620] = 0; 
  adj[3621] = 0; 
  adj[3622] = 0; 
  adj[3623] = 0; 
  adj[3624] = 0; 
  adj[3625] = 0; 
  adj[3626] = 0; 
  adj[3627] = 0; 
  adj[3628] = 0; 
  adj[3629] = 0; 
  adj[3630] = 0; 
  adj[3631] = 0; 
  adj[3632] = 0; 
  adj[3633] = 0; 
  adj[3634] = 0; 
  adj[3635] = 0; 
  adj[3636] = 0; 
  adj[3637] = 0; 
  adj[3638] = 0; 
  adj[3639] = 1; 
  adj[3640] = 0; 
  adj[3641] = 1; 
  adj[3642] = 0; 
  adj[3643] = 0; 
  adj[3644] = 0; 
  adj[3645] = 0; 
  adj[3646] = 0; 
  adj[3647] = 0; 
  adj[3648] = 0; 
  adj[3649] = 0; 
  adj[3650] = 0; 
  adj[3651] = 0; 
  adj[3652] = 0; 
  adj[3653] = 0; 
  adj[3654] = 0; 
  adj[3655] = 0; 
  adj[3656] = 0; 
  adj[3657] = 0; 
  adj[3658] = 0; 
  adj[3659] = 0; 
  adj[3660] = 0; 
  adj[3661] = 0; 
  adj[3662] = 0; 
  adj[3663] = 0; 
  adj[3664] = 0; 
  adj[3665] = 0; 
  adj[3666] = 0; 
  adj[3667] = 0; 
  adj[3668] = 0; 
  adj[3669] = 0; 
  adj[3670] = 0; 
  adj[3671] = 0; 
  adj[3672] = 0; 
  adj[3673] = 0; 
  adj[3674] = 0; 
  adj[3675] = 0; 
  adj[3676] = 0; 
  adj[3677] = 0; 
  adj[3678] = 0; 
  adj[3679] = 0; 
  adj[3680] = 0; 
  adj[3681] = 0; 
  adj[3682] = 0; 
  adj[3683] = 0; 
  adj[3684] = 0; 
  adj[3685] = 0; 
  adj[3686] = 0; 
  adj[3687] = 0; 
  adj[3688] = 0; 
  adj[3689] = 0; 
  adj[3690] = 0; 
  adj[3691] = 0; 
  adj[3692] = 0; 
  adj[3693] = 0; 
  adj[3694] = 0; 
  adj[3695] = 0; 
  adj[3696] = 0; 
  adj[3697] = 0; 
  adj[3698] = 0; 
  adj[3699] = 0; 
  adj[3700] = 0; 
  adj[3701] = 0; 
  adj[3702] = 0; 
  adj[3703] = 0; 
  adj[3704] = 1; 
  adj[3705] = 0; 
  adj[3706] = 1; 
  adj[3707] = 0; 
  adj[3708] = 0; 
  adj[3709] = 0; 
  adj[3710] = 0; 
  adj[3711] = 0; 
  adj[3712] = 0; 
  adj[3713] = 0; 
  adj[3714] = 0; 
  adj[3715] = 0; 
  adj[3716] = 0; 
  adj[3717] = 0; 
  adj[3718] = 0; 
  adj[3719] = 0; 
  adj[3720] = 0; 
  adj[3721] = 0; 
  adj[3722] = 0; 
  adj[3723] = 0; 
  adj[3724] = 0; 
  adj[3725] = 0; 
  adj[3726] = 0; 
  adj[3727] = 0; 
  adj[3728] = 0; 
  adj[3729] = 0; 
  adj[3730] = 0; 
  adj[3731] = 0; 
  adj[3732] = 0; 
  adj[3733] = 0; 
  adj[3734] = 0; 
  adj[3735] = 0; 
  adj[3736] = 0; 
  adj[3737] = 0; 
  adj[3738] = 0; 
  adj[3739] = 0; 
  adj[3740] = 0; 
  adj[3741] = 0; 
  adj[3742] = 0; 
  adj[3743] = 0; 
  adj[3744] = 0; 
  adj[3745] = 0; 
  adj[3746] = 0; 
  adj[3747] = 0; 
  adj[3748] = 0; 
  adj[3749] = 0; 
  adj[3750] = 0; 
  adj[3751] = 0; 
  adj[3752] = 0; 
  adj[3753] = 0; 
  adj[3754] = 0; 
  adj[3755] = 0; 
  adj[3756] = 0; 
  adj[3757] = 0; 
  adj[3758] = 0; 
  adj[3759] = 0; 
  adj[3760] = 0; 
  adj[3761] = 0; 
  adj[3762] = 0; 
  adj[3763] = 0; 
  adj[3764] = 0; 
  adj[3765] = 0; 
  adj[3766] = 0; 
  adj[3767] = 0; 
  adj[3768] = 0; 
  adj[3769] = 1; 
  adj[3770] = 0; 
  adj[3771] = 1; 
  adj[3772] = 0; 
  adj[3773] = 0; 
  adj[3774] = 0; 
  adj[3775] = 0; 
  adj[3776] = 0; 
  adj[3777] = 0; 
  adj[3778] = 0; 
  adj[3779] = 0; 
  adj[3780] = 0; 
  adj[3781] = 0; 
  adj[3782] = 0; 
  adj[3783] = 0; 
  adj[3784] = 0; 
  adj[3785] = 0; 
  adj[3786] = 0; 
  adj[3787] = 0; 
  adj[3788] = 0; 
  adj[3789] = 0; 
  adj[3790] = 0; 
  adj[3791] = 0; 
  adj[3792] = 0; 
  adj[3793] = 0; 
  adj[3794] = 0; 
  adj[3795] = 0; 
  adj[3796] = 0; 
  adj[3797] = 0; 
  adj[3798] = 0; 
  adj[3799] = 0; 
  adj[3800] = 0; 
  adj[3801] = 0; 
  adj[3802] = 0; 
  adj[3803] = 0; 
  adj[3804] = 0; 
  adj[3805] = 0; 
  adj[3806] = 0; 
  adj[3807] = 0; 
  adj[3808] = 0; 
  adj[3809] = 0; 
  adj[3810] = 0; 
  adj[3811] = 0; 
  adj[3812] = 0; 
  adj[3813] = 0; 
  adj[3814] = 0; 
  adj[3815] = 0; 
  adj[3816] = 0; 
  adj[3817] = 0; 
  adj[3818] = 0; 
  adj[3819] = 0; 
  adj[3820] = 0; 
  adj[3821] = 0; 
  adj[3822] = 0; 
  adj[3823] = 0; 
  adj[3824] = 0; 
  adj[3825] = 0; 
  adj[3826] = 0; 
  adj[3827] = 0; 
  adj[3828] = 0; 
  adj[3829] = 0; 
  adj[3830] = 0; 
  adj[3831] = 0; 
  adj[3832] = 0; 
  adj[3833] = 0; 
  adj[3834] = 1; 
  adj[3835] = 0; 
  adj[3836] = 1; 
  adj[3837] = 0; 
  adj[3838] = 0; 
  adj[3839] = 0; 
  adj[3840] = 0; 
  adj[3841] = 0; 
  adj[3842] = 0; 
  adj[3843] = 0; 
  adj[3844] = 0; 
  adj[3845] = 0; 
  adj[3846] = 0; 
  adj[3847] = 0; 
  adj[3848] = 0; 
  adj[3849] = 0; 
  adj[3850] = 0; 
  adj[3851] = 0; 
  adj[3852] = 0; 
  adj[3853] = 0; 
  adj[3854] = 0; 
  adj[3855] = 0; 
  adj[3856] = 0; 
  adj[3857] = 0; 
  adj[3858] = 0; 
  adj[3859] = 0; 
  adj[3860] = 0; 
  adj[3861] = 0; 
  adj[3862] = 0; 
  adj[3863] = 0; 
  adj[3864] = 0; 
  adj[3865] = 0; 
  adj[3866] = 0; 
  adj[3867] = 0; 
  adj[3868] = 0; 
  adj[3869] = 0; 
  adj[3870] = 0; 
  adj[3871] = 0; 
  adj[3872] = 0; 
  adj[3873] = 0; 
  adj[3874] = 0; 
  adj[3875] = 0; 
  adj[3876] = 0; 
  adj[3877] = 0; 
  adj[3878] = 0; 
  adj[3879] = 0; 
  adj[3880] = 0; 
  adj[3881] = 0; 
  adj[3882] = 0; 
  adj[3883] = 0; 
  adj[3884] = 0; 
  adj[3885] = 0; 
  adj[3886] = 0; 
  adj[3887] = 0; 
  adj[3888] = 0; 
  adj[3889] = 0; 
  adj[3890] = 0; 
  adj[3891] = 0; 
  adj[3892] = 0; 
  adj[3893] = 0; 
  adj[3894] = 0; 
  adj[3895] = 0; 
  adj[3896] = 0; 
  adj[3897] = 0; 
  adj[3898] = 0; 
  adj[3899] = 1; 
  adj[3900] = 0; 
  adj[3901] = 1; 
  adj[3902] = 0; 
  adj[3903] = 0; 
  adj[3904] = 0; 
  adj[3905] = 0; 
  adj[3906] = 0; 
  adj[3907] = 0; 
  adj[3908] = 0; 
  adj[3909] = 0; 
  adj[3910] = 0; 
  adj[3911] = 0; 
  adj[3912] = 0; 
  adj[3913] = 0; 
  adj[3914] = 0; 
  adj[3915] = 0; 
  adj[3916] = 0; 
  adj[3917] = 0; 
  adj[3918] = 0; 
  adj[3919] = 0; 
  adj[3920] = 0; 
  adj[3921] = 0; 
  adj[3922] = 0; 
  adj[3923] = 0; 
  adj[3924] = 0; 
  adj[3925] = 0; 
  adj[3926] = 0; 
  adj[3927] = 0; 
  adj[3928] = 0; 
  adj[3929] = 0; 
  adj[3930] = 0; 
  adj[3931] = 0; 
  adj[3932] = 0; 
  adj[3933] = 0; 
  adj[3934] = 0; 
  adj[3935] = 0; 
  adj[3936] = 0; 
  adj[3937] = 0; 
  adj[3938] = 0; 
  adj[3939] = 0; 
  adj[3940] = 0; 
  adj[3941] = 0; 
  adj[3942] = 0; 
  adj[3943] = 0; 
  adj[3944] = 0; 
  adj[3945] = 0; 
  adj[3946] = 0; 
  adj[3947] = 0; 
  adj[3948] = 0; 
  adj[3949] = 0; 
  adj[3950] = 0; 
  adj[3951] = 0; 
  adj[3952] = 0; 
  adj[3953] = 0; 
  adj[3954] = 0; 
  adj[3955] = 0; 
  adj[3956] = 0; 
  adj[3957] = 0; 
  adj[3958] = 0; 
  adj[3959] = 0; 
  adj[3960] = 0; 
  adj[3961] = 0; 
  adj[3962] = 0; 
  adj[3963] = 0; 
  adj[3964] = 1; 
  adj[3965] = 0; 
  adj[3966] = 1; 
  adj[3967] = 0; 
  adj[3968] = 0; 
  adj[3969] = 0; 
  adj[3970] = 0; 
  adj[3971] = 0; 
  adj[3972] = 0; 
  adj[3973] = 0; 
  adj[3974] = 0; 
  adj[3975] = 0; 
  adj[3976] = 0; 
  adj[3977] = 0; 
  adj[3978] = 0; 
  adj[3979] = 0; 
  adj[3980] = 0; 
  adj[3981] = 0; 
  adj[3982] = 0; 
  adj[3983] = 0; 
  adj[3984] = 0; 
  adj[3985] = 0; 
  adj[3986] = 0; 
  adj[3987] = 0; 
  adj[3988] = 0; 
  adj[3989] = 0; 
  adj[3990] = 0; 
  adj[3991] = 0; 
  adj[3992] = 0; 
  adj[3993] = 0; 
  adj[3994] = 0; 
  adj[3995] = 0; 
  adj[3996] = 0; 
  adj[3997] = 0; 
  adj[3998] = 0; 
  adj[3999] = 0; 
  adj[4000] = 0; 
  adj[4001] = 0; 
  adj[4002] = 0; 
  adj[4003] = 0; 
  adj[4004] = 0; 
  adj[4005] = 0; 
  adj[4006] = 0; 
  adj[4007] = 0; 
  adj[4008] = 0; 
  adj[4009] = 0; 
  adj[4010] = 0; 
  adj[4011] = 0; 
  adj[4012] = 0; 
  adj[4013] = 0; 
  adj[4014] = 0; 
  adj[4015] = 0; 
  adj[4016] = 0; 
  adj[4017] = 0; 
  adj[4018] = 0; 
  adj[4019] = 0; 
  adj[4020] = 0; 
  adj[4021] = 0; 
  adj[4022] = 0; 
  adj[4023] = 0; 
  adj[4024] = 0; 
  adj[4025] = 0; 
  adj[4026] = 0; 
  adj[4027] = 0; 
  adj[4028] = 0; 
  adj[4029] = 1; 
  adj[4030] = 0; 
  adj[4031] = 1; 
  adj[4032] = 1; 
  adj[4033] = 0; 
  adj[4034] = 0; 
  adj[4035] = 0; 
  adj[4036] = 0; 
  adj[4037] = 0; 
  adj[4038] = 0; 
  adj[4039] = 0; 
  adj[4040] = 0; 
  adj[4041] = 0; 
  adj[4042] = 0; 
  adj[4043] = 0; 
  adj[4044] = 1; 
  adj[4045] = 0; 
  adj[4046] = 0; 
  adj[4047] = 0; 
  adj[4048] = 0; 
  adj[4049] = 0; 
  adj[4050] = 0; 
  adj[4051] = 0; 
  adj[4052] = 0; 
  adj[4053] = 0; 
  adj[4054] = 0; 
  adj[4055] = 0; 
  adj[4056] = 0; 
  adj[4057] = 0; 
  adj[4058] = 0; 
  adj[4059] = 0; 
  adj[4060] = 0; 
  adj[4061] = 0; 
  adj[4062] = 0; 
  adj[4063] = 0; 
  adj[4064] = 0; 
  adj[4065] = 0; 
  adj[4066] = 0; 
  adj[4067] = 0; 
  adj[4068] = 0; 
  adj[4069] = 0; 
  adj[4070] = 0; 
  adj[4071] = 0; 
  adj[4072] = 0; 
  adj[4073] = 0; 
  adj[4074] = 0; 
  adj[4075] = 0; 
  adj[4076] = 0; 
  adj[4077] = 0; 
  adj[4078] = 0; 
  adj[4079] = 0; 
  adj[4080] = 0; 
  adj[4081] = 0; 
  adj[4082] = 0; 
  adj[4083] = 0; 
  adj[4084] = 0; 
  adj[4085] = 0; 
  adj[4086] = 0; 
  adj[4087] = 0; 
  adj[4088] = 0; 
  adj[4089] = 0; 
  adj[4090] = 0; 
  adj[4091] = 0; 
  adj[4092] = 0; 
  adj[4093] = 0; 
  adj[4094] = 1; 
  adj[4095] = 0; 
  nodeWeight[1*WIDTH-1:0*WIDTH] =  16'h8000; 
  nodeWeight[2*WIDTH-1:1*WIDTH] =  16'h8000; 
  nodeWeight[3*WIDTH-1:2*WIDTH] =  16'h8000; 
  nodeWeight[4*WIDTH-1:3*WIDTH] =  16'h8000; 
  nodeWeight[5*WIDTH-1:4*WIDTH] =  16'h8000; 
  nodeWeight[6*WIDTH-1:5*WIDTH] =  16'h8000; 
  nodeWeight[7*WIDTH-1:6*WIDTH] =  16'h8000; 
  nodeWeight[8*WIDTH-1:7*WIDTH] =  16'h8000; 
  nodeWeight[9*WIDTH-1:8*WIDTH] =  16'h8000; 
  nodeWeight[10*WIDTH-1:9*WIDTH] =  16'h8000; 
  nodeWeight[11*WIDTH-1:10*WIDTH] =  16'h8000; 
  nodeWeight[12*WIDTH-1:11*WIDTH] =  16'h8000; 
  nodeWeight[13*WIDTH-1:12*WIDTH] =  16'h5555; 
  nodeWeight[14*WIDTH-1:13*WIDTH] =  16'h8000; 
  nodeWeight[15*WIDTH-1:14*WIDTH] =  16'h8000; 
  nodeWeight[16*WIDTH-1:15*WIDTH] =  16'h8000; 
  nodeWeight[17*WIDTH-1:16*WIDTH] =  16'h8000; 
  nodeWeight[18*WIDTH-1:17*WIDTH] =  16'h5555; 
  nodeWeight[19*WIDTH-1:18*WIDTH] =  16'h8000; 
  nodeWeight[20*WIDTH-1:19*WIDTH] =  16'h8000; 
  nodeWeight[21*WIDTH-1:20*WIDTH] =  16'h8000; 
  nodeWeight[22*WIDTH-1:21*WIDTH] =  16'h5555; 
  nodeWeight[23*WIDTH-1:22*WIDTH] =  16'h8000; 
  nodeWeight[24*WIDTH-1:23*WIDTH] =  16'h8000; 
  nodeWeight[25*WIDTH-1:24*WIDTH] =  16'h8000; 
  nodeWeight[26*WIDTH-1:25*WIDTH] =  16'h8000; 
  nodeWeight[27*WIDTH-1:26*WIDTH] =  16'h8000; 
  nodeWeight[28*WIDTH-1:27*WIDTH] =  16'h4000; 
  nodeWeight[29*WIDTH-1:28*WIDTH] =  16'h8000; 
  nodeWeight[30*WIDTH-1:29*WIDTH] =  16'h8000; 
  nodeWeight[31*WIDTH-1:30*WIDTH] =  16'h8000; 
  nodeWeight[32*WIDTH-1:31*WIDTH] =  16'h8000; 
  nodeWeight[33*WIDTH-1:32*WIDTH] =  16'h8000; 
  nodeWeight[34*WIDTH-1:33*WIDTH] =  16'h8000; 
  nodeWeight[35*WIDTH-1:34*WIDTH] =  16'h8000; 
  nodeWeight[36*WIDTH-1:35*WIDTH] =  16'h8000; 
  nodeWeight[37*WIDTH-1:36*WIDTH] =  16'h8000; 
  nodeWeight[38*WIDTH-1:37*WIDTH] =  16'h8000; 
  nodeWeight[39*WIDTH-1:38*WIDTH] =  16'h8000; 
  nodeWeight[40*WIDTH-1:39*WIDTH] =  16'h5555; 
  nodeWeight[41*WIDTH-1:40*WIDTH] =  16'h8000; 
  nodeWeight[42*WIDTH-1:41*WIDTH] =  16'h8000; 
  nodeWeight[43*WIDTH-1:42*WIDTH] =  16'h8000; 
  nodeWeight[44*WIDTH-1:43*WIDTH] =  16'h8000; 
  nodeWeight[45*WIDTH-1:44*WIDTH] =  16'h8000; 
  nodeWeight[46*WIDTH-1:45*WIDTH] =  16'h8000; 
  nodeWeight[47*WIDTH-1:46*WIDTH] =  16'h8000; 
  nodeWeight[48*WIDTH-1:47*WIDTH] =  16'h8000; 
  nodeWeight[49*WIDTH-1:48*WIDTH] =  16'h8000; 
  nodeWeight[50*WIDTH-1:49*WIDTH] =  16'h8000; 
  nodeWeight[51*WIDTH-1:50*WIDTH] =  16'h8000; 
  nodeWeight[52*WIDTH-1:51*WIDTH] =  16'h8000; 
  nodeWeight[53*WIDTH-1:52*WIDTH] =  16'h5555; 
  nodeWeight[54*WIDTH-1:53*WIDTH] =  16'h8000; 
  nodeWeight[55*WIDTH-1:54*WIDTH] =  16'h8000; 
  nodeWeight[56*WIDTH-1:55*WIDTH] =  16'h8000; 
  nodeWeight[57*WIDTH-1:56*WIDTH] =  16'h8000; 
  nodeWeight[58*WIDTH-1:57*WIDTH] =  16'h8000; 
  nodeWeight[59*WIDTH-1:58*WIDTH] =  16'h8000; 
  nodeWeight[60*WIDTH-1:59*WIDTH] =  16'h8000; 
  nodeWeight[61*WIDTH-1:60*WIDTH] =  16'h8000; 
  nodeWeight[62*WIDTH-1:61*WIDTH] =  16'h8000; 
  nodeWeight[63*WIDTH-1:62*WIDTH] =  16'h8000; 
  nodeWeight[64*WIDTH-1:63*WIDTH] =  16'h5555; 

	#2 reset = 1'b0;
end

endmodule
